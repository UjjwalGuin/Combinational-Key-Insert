
module b15 ( BE_n, Address, W_R_n, D_C_n, M_IO_n, ADS_n, Datai, Datao, CK, 
        NA_n, BS16_n, READY_n, HOLD, reset );
  output [3:0] BE_n;
  output [29:0] Address;
  input [31:0] Datai;
  output [31:0] Datao;
  input CK, NA_n, BS16_n, READY_n, HOLD, reset;
  output W_R_n, D_C_n, M_IO_n, ADS_n;
  wire   n730, n731, n732, n755, n789, n790, n791, n792, n801, n803, n805,
         n807, n809, n811, n813, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n965, n973, n974,
         n975, n976, n979, n4488, n4489, n4490, n4491, n4492, n4493, n4494,
         n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504,
         n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514,
         n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524,
         n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534,
         n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544,
         n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554,
         n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564,
         n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574,
         n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584,
         n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594,
         n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604,
         n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614,
         n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624,
         n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634,
         n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644,
         n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654,
         n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664,
         n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674,
         n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684,
         n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694,
         n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704,
         n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714,
         n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724,
         n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734,
         n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744,
         n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754,
         n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764,
         n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774,
         n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784,
         n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794,
         n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804,
         n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814,
         n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824,
         n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834,
         n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844,
         n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854,
         n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864,
         n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874,
         n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884,
         n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894,
         n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905,
         n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915,
         n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925,
         n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935,
         n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945,
         n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955,
         n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965,
         n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975,
         n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985,
         n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995,
         n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005,
         n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015,
         n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025,
         n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035,
         n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045,
         n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055,
         n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065,
         n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075,
         n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085,
         n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095,
         n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105,
         n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115,
         n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125,
         n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135,
         n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145,
         n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155,
         n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165,
         n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175,
         n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185,
         n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195,
         n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205,
         n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215,
         n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225,
         n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235,
         n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245,
         n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255,
         n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265,
         n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275,
         n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285,
         n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295,
         n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305,
         n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315,
         n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325,
         n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335,
         n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345,
         n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355,
         n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365,
         n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375,
         n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385,
         n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395,
         n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405,
         n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415,
         n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425,
         n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435,
         n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445,
         n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455,
         n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465,
         n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475,
         n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485,
         n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495,
         n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505,
         n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515,
         n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525,
         n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535,
         n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545,
         n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555,
         n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565,
         n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575,
         n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585,
         n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595,
         n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605,
         n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615,
         n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625,
         n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635,
         n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645,
         n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655,
         n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665,
         n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675,
         n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685,
         n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695,
         n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705,
         n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715,
         n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725,
         n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735,
         n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745,
         n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755,
         n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765,
         n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775,
         n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785,
         n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795,
         n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805,
         n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815,
         n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825,
         n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835,
         n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845,
         n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855,
         n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865,
         n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875,
         n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885,
         n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895,
         n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905,
         n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915,
         n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925,
         n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935,
         n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945,
         n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955,
         n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965,
         n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975,
         n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985,
         n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995,
         n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005,
         n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015,
         n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025,
         n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035,
         n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045,
         n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055,
         n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065,
         n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075,
         n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085,
         n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095,
         n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105,
         n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115,
         n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125,
         n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135,
         n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145,
         n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155,
         n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165,
         n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175,
         n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185,
         n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195,
         n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205,
         n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215,
         n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225,
         n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235,
         n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245,
         n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255,
         n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265,
         n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275,
         n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285,
         n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295,
         n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305,
         n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315,
         n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325,
         n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335,
         n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345,
         n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355,
         n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365,
         n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375,
         n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385,
         n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395,
         n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405,
         n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415,
         n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425,
         n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435,
         n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445,
         n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455,
         n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465,
         n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475,
         n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485,
         n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495,
         n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505,
         n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515,
         n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525,
         n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535,
         n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545,
         n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555,
         n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565,
         n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575,
         n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585,
         n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595,
         n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605,
         n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615,
         n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625,
         n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635,
         n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645,
         n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655,
         n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665,
         n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675,
         n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685,
         n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695,
         n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705,
         n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715,
         n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725,
         n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735,
         n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745,
         n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755,
         n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765,
         n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775,
         n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785,
         n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795,
         n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805,
         n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815,
         n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825,
         n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835,
         n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845,
         n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855,
         n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865,
         n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875,
         n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885,
         n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895,
         n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905,
         n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915,
         n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925,
         n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935,
         n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945,
         n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955,
         n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965,
         n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975,
         n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985,
         n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995,
         n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005,
         n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015,
         n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025,
         n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035,
         n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045,
         n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055,
         n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065,
         n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075,
         n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085,
         n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095,
         n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105,
         n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115,
         n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125,
         n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135,
         n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145,
         n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155,
         n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165,
         n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175,
         n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185,
         n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195,
         n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205,
         n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215,
         n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225,
         n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235,
         n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245,
         n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255,
         n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265,
         n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275,
         n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285,
         n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295,
         n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305,
         n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315,
         n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325,
         n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335,
         n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345,
         n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355,
         n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365,
         n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375,
         n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385,
         n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395,
         n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405,
         n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415,
         n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425,
         n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435,
         n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445,
         n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455,
         n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465,
         n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475,
         n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485,
         n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495,
         n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505,
         n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515,
         n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525,
         n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535,
         n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545,
         n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555,
         n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565,
         n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575,
         n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585,
         n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595,
         n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605,
         n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615,
         n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625,
         n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635,
         n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645,
         n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655,
         n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665,
         n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675,
         n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685,
         n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695,
         n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705,
         n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715,
         n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725,
         n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735,
         n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745,
         n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755,
         n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765,
         n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775,
         n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785,
         n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795,
         n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805,
         n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815,
         n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825,
         n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835,
         n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845,
         n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855,
         n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865,
         n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875,
         n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885,
         n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895,
         n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905,
         n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915,
         n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925,
         n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935,
         n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945,
         n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955,
         n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965,
         n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975,
         n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985,
         n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995,
         n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005,
         n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015,
         n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025,
         n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035,
         n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045,
         n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055,
         n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065,
         n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075,
         n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085,
         n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095,
         n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105,
         n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115,
         n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125,
         n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135,
         n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145,
         n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155,
         n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165,
         n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175,
         n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185,
         n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195,
         n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205,
         n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215,
         n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225,
         n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235,
         n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245,
         n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255,
         n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265,
         n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275,
         n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285,
         n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295,
         n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305,
         n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315,
         n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325,
         n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335,
         n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345,
         n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355,
         n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365,
         n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375,
         n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385,
         n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395,
         n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405,
         n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415,
         n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425,
         n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435,
         n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445,
         n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455,
         n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465,
         n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475,
         n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485,
         n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495,
         n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505,
         n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515,
         n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525,
         n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535,
         n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545,
         n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555,
         n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565,
         n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575,
         n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585,
         n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595,
         n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605,
         n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615,
         n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625,
         n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635,
         n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645,
         n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655,
         n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665,
         n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675,
         n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685,
         n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695,
         n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705,
         n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715,
         n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725,
         n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735,
         n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745,
         n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755,
         n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765,
         n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775,
         n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785,
         n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795,
         n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805,
         n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815,
         n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825,
         n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835,
         n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845,
         n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855,
         n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865,
         n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875,
         n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885,
         n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895,
         n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905,
         n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915,
         n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925,
         n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935,
         n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945,
         n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955,
         n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965,
         n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975,
         n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985,
         n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995,
         n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005,
         n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015,
         n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025,
         n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035,
         n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045,
         n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055,
         n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065,
         n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075,
         n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085,
         n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095,
         n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105,
         n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115,
         n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125,
         n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135,
         n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145,
         n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155,
         n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165,
         n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175,
         n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185,
         n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195,
         n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205,
         n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215,
         n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225,
         n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235,
         n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245,
         n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255,
         n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265,
         n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275,
         n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285,
         n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295,
         n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305,
         n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315,
         n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325,
         n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335,
         n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345,
         n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355,
         n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365,
         n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375,
         n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385,
         n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395,
         n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405,
         n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415,
         n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425,
         n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435,
         n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445,
         n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455,
         n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465,
         n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475,
         n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485,
         n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495,
         n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505,
         n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515,
         n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525,
         n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535,
         n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545,
         n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555,
         n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565,
         n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575,
         n9576, n9577, n9578, n9579, n9580, n9581;
  wire   [31:0] rEIP;
  wire   [14:0] uWord;
  assign Datao[31] = 1'b0;
  //add;

  //gate;
  DFFARX1_RVT RequestPending_reg ( .D(n4904), .CLK(CK), .RSTB(n5250), .Q(n4989), .QN(n979) );
  DFFARX1_RVT State_reg_2_ ( .D(n4903), .CLK(CK), .RSTB(n5250), .Q(n4913), 
        .QN(n730) );
  DFFARX1_RVT State_reg_1_ ( .D(n4901), .CLK(CK), .RSTB(n5250), .Q(n4962), 
        .QN(n731) );
  DFFARX1_RVT State_reg_0_ ( .D(n4902), .CLK(CK), .RSTB(n5250), .Q(n4929), 
        .QN(n732) );
  DFFARX1_RVT ADS_n_reg ( .D(n4900), .CLK(CK), .RSTB(n5250), .Q(ADS_n) );
  DFFARX1_RVT StateBS16_reg ( .D(n4899), .CLK(CK), .RSTB(n5250), .Q(n4967), 
        .QN(n755) );
  DFFARX1_RVT PhyAddrPointer_reg_31_ ( .D(n4527), .CLK(CK), .RSTB(n5219), .Q(
        n5086) );
  DFFARX1_RVT rEIP_reg_31_ ( .D(n4589), .CLK(CK), .RSTB(n5219), .Q(rEIP[31])
         );
  DFFARX1_RVT InstAddrPointer_reg_31_ ( .D(n4896), .CLK(CK), .RSTB(n5247), 
        .QN(n9567) );
  DFFARX1_RVT InstQueueRd_Addr_reg_1_ ( .D(n4758), .CLK(CK), .RSTB(n5247), .Q(
        n4927), .QN(n938) );
  DFFARX1_RVT EBX_reg_31_ ( .D(n4621), .CLK(CK), .RSTB(n5220), .Q(n4958) );
  DFFARX1_RVT rEIP_reg_30_ ( .D(n4590), .CLK(CK), .RSTB(n5219), .Q(rEIP[30])
         );
  DFFARX1_RVT InstAddrPointer_reg_30_ ( .D(n4752), .CLK(CK), .RSTB(n5247), 
        .QN(n9568) );
  DFFARX1_RVT PhyAddrPointer_reg_0_ ( .D(n4558), .CLK(CK), .RSTB(n5235), .Q(
        n5055) );
  DFFARX1_RVT rEIP_reg_0_ ( .D(n4620), .CLK(CK), .RSTB(n5249), .Q(rEIP[0]) );
  DFFARX1_RVT InstAddrPointer_reg_0_ ( .D(n4753), .CLK(CK), .RSTB(n5249), .Q(
        n4931), .QN(n976) );
  DFFARX1_RVT InstQueueRd_Addr_reg_0_ ( .D(n4761), .CLK(CK), .RSTB(n5247), .Q(
        n4908), .QN(n939) );
  DFFARX1_RVT State2_reg_1_ ( .D(n4755), .CLK(CK), .RSTB(n5246), .Q(n4910), 
        .QN(n791) );
  DFFARX1_RVT State2_reg_0_ ( .D(n4757), .CLK(CK), .RSTB(n5249), .Q(n4969), 
        .QN(n792) );
  DFFARX1_RVT State2_reg_3_ ( .D(n4893), .CLK(CK), .RSTB(n5246), .Q(n4925), 
        .QN(n789) );
  DFFARX1_RVT State2_reg_2_ ( .D(n4756), .CLK(CK), .RSTB(n5246), .Q(n4905), 
        .QN(n790) );
  DFFARX1_RVT CodeFetch_reg ( .D(n4717), .CLK(CK), .RSTB(n5239), .Q(n5195), 
        .QN(n9511) );
  DFFARX1_RVT D_C_n_reg ( .D(n4716), .CLK(CK), .RSTB(n5239), .Q(D_C_n) );
  DFFARX1_RVT Flush_reg ( .D(n4754), .CLK(CK), .RSTB(n5246), .Q(n5110), .QN(
        n9561) );
  DFFARX1_RVT InstQueueWr_Addr_reg_0_ ( .D(n4891), .CLK(CK), .RSTB(n5247), .Q(
        n4928), .QN(n975) );
  DFFARX1_RVT InstQueueWr_Addr_reg_1_ ( .D(n4892), .CLK(CK), .RSTB(n5247), .Q(
        n4909), .QN(n974) );
  DFFARX1_RVT InstQueueWr_Addr_reg_2_ ( .D(n4890), .CLK(CK), .RSTB(n5247), .Q(
        n4907), .QN(n973) );
  DFFARX1_RVT InstQueueWr_Addr_reg_3_ ( .D(n4889), .CLK(CK), .RSTB(n5247), .Q(
        n4930), .QN(n965) );
  DFFARX1_RVT InstQueue_reg_14__7_ ( .D(n4769), .CLK(CK), .RSTB(n5244), .Q(
        n5048), .QN(n816) );
  DFFARX1_RVT MemoryFetch_reg ( .D(n4719), .CLK(CK), .RSTB(n5239), .Q(n5173)
         );
  DFFARX1_RVT M_IO_n_reg ( .D(n4718), .CLK(CK), .RSTB(n5239), .Q(M_IO_n) );
  DFFARX1_RVT InstQueueRd_Addr_reg_2_ ( .D(n4759), .CLK(CK), .RSTB(n5249), .Q(
        n4926), .QN(n937) );
  DFFARX1_RVT InstQueue_reg_0__2_ ( .D(n4886), .CLK(CK), .RSTB(n5246), .Q(
        n5131), .QN(n933) );
  DFFARX1_RVT InstQueue_reg_1__2_ ( .D(n4878), .CLK(CK), .RSTB(n5236), .Q(
        n5130), .QN(n925) );
  DFFARX1_RVT InstQueue_reg_2__2_ ( .D(n4870), .CLK(CK), .RSTB(n5236), .Q(
        n5142), .QN(n917) );
  DFFARX1_RVT InstQueue_reg_3__2_ ( .D(n4862), .CLK(CK), .RSTB(n5236), .Q(
        n5146), .QN(n909) );
  DFFARX1_RVT InstQueue_reg_4__2_ ( .D(n4854), .CLK(CK), .RSTB(n5237), .Q(
        n5144), .QN(n901) );
  DFFARX1_RVT InstQueue_reg_5__2_ ( .D(n4846), .CLK(CK), .RSTB(n5237), .Q(
        n5011), .QN(n893) );
  DFFARX1_RVT InstQueue_reg_6__2_ ( .D(n4838), .CLK(CK), .RSTB(n5237), .Q(
        n5014), .QN(n885) );
  DFFARX1_RVT InstQueue_reg_7__2_ ( .D(n4830), .CLK(CK), .RSTB(n5237), .Q(
        n5108), .QN(n877) );
  DFFARX1_RVT InstQueue_reg_8__2_ ( .D(n4822), .CLK(CK), .RSTB(n5237), .Q(
        n5145), .QN(n869) );
  DFFARX1_RVT InstQueue_reg_9__2_ ( .D(n4814), .CLK(CK), .RSTB(n5237), .Q(
        n5012), .QN(n861) );
  DFFARX1_RVT InstQueue_reg_10__2_ ( .D(n4806), .CLK(CK), .RSTB(n5237), .Q(
        n5013), .QN(n853) );
  DFFARX1_RVT InstQueue_reg_11__2_ ( .D(n4798), .CLK(CK), .RSTB(n5237), .Q(
        n5015), .QN(n845) );
  DFFARX1_RVT InstQueue_reg_12__2_ ( .D(n4790), .CLK(CK), .RSTB(n5237), .Q(
        n5143), .QN(n837) );
  DFFARX1_RVT InstQueue_reg_13__2_ ( .D(n4782), .CLK(CK), .RSTB(n5237), .Q(
        n5010), .QN(n829) );
  DFFARX1_RVT InstQueue_reg_14__2_ ( .D(n4774), .CLK(CK), .RSTB(n5237), .Q(
        n5113), .QN(n821) );
  DFFARX1_RVT InstQueue_reg_15__2_ ( .D(n4766), .CLK(CK), .RSTB(n5237), .QN(
        n811) );
  DFFARX1_RVT InstQueue_reg_15__3_ ( .D(n4765), .CLK(CK), .RSTB(n5239), .QN(
        n809) );
  DFFARX1_RVT InstQueue_reg_14__3_ ( .D(n4773), .CLK(CK), .RSTB(n5239), .Q(
        n5114), .QN(n820) );
  DFFARX1_RVT InstQueue_reg_13__3_ ( .D(n4781), .CLK(CK), .RSTB(n5239), .Q(
        n5016), .QN(n828) );
  DFFARX1_RVT InstQueue_reg_12__3_ ( .D(n4789), .CLK(CK), .RSTB(n5238), .Q(
        n5148), .QN(n836) );
  DFFARX1_RVT InstQueue_reg_11__3_ ( .D(n4797), .CLK(CK), .RSTB(n5238), .Q(
        n5021), .QN(n844) );
  DFFARX1_RVT InstQueue_reg_10__3_ ( .D(n4805), .CLK(CK), .RSTB(n5238), .Q(
        n5019), .QN(n852) );
  DFFARX1_RVT InstQueue_reg_9__3_ ( .D(n4813), .CLK(CK), .RSTB(n5238), .Q(
        n5018), .QN(n860) );
  DFFARX1_RVT InstQueue_reg_8__3_ ( .D(n4821), .CLK(CK), .RSTB(n5238), .Q(
        n5150), .QN(n868) );
  DFFARX1_RVT InstQueue_reg_7__3_ ( .D(n4829), .CLK(CK), .RSTB(n5238), .Q(
        n5022), .QN(n876) );
  DFFARX1_RVT InstQueue_reg_6__3_ ( .D(n4837), .CLK(CK), .RSTB(n5238), .Q(
        n5020), .QN(n884) );
  DFFARX1_RVT InstQueue_reg_5__3_ ( .D(n4845), .CLK(CK), .RSTB(n5238), .Q(
        n5017), .QN(n892) );
  DFFARX1_RVT InstQueue_reg_4__3_ ( .D(n4853), .CLK(CK), .RSTB(n5238), .Q(
        n5149), .QN(n900) );
  DFFARX1_RVT InstQueue_reg_3__3_ ( .D(n4861), .CLK(CK), .RSTB(n5238), .Q(
        n5151), .QN(n908) );
  DFFARX1_RVT InstQueue_reg_2__3_ ( .D(n4869), .CLK(CK), .RSTB(n5238), .Q(
        n5147), .QN(n916) );
  DFFARX1_RVT InstQueue_reg_1__3_ ( .D(n4877), .CLK(CK), .RSTB(n5238), .Q(
        n5124), .QN(n924) );
  DFFARX1_RVT InstQueue_reg_0__3_ ( .D(n4885), .CLK(CK), .RSTB(n5246), .Q(
        n5119), .QN(n932) );
  DFFARX1_RVT InstQueue_reg_15__1_ ( .D(n4767), .CLK(CK), .RSTB(n5240), .QN(
        n813) );
  DFFARX1_RVT InstQueue_reg_14__1_ ( .D(n4775), .CLK(CK), .RSTB(n5240), .Q(
        n5112), .QN(n822) );
  DFFARX1_RVT InstQueue_reg_13__1_ ( .D(n4783), .CLK(CK), .RSTB(n5240), .Q(
        n5003), .QN(n830) );
  DFFARX1_RVT InstQueue_reg_12__1_ ( .D(n4791), .CLK(CK), .RSTB(n5240), .Q(
        n5138), .QN(n838) );
  DFFARX1_RVT InstQueue_reg_11__1_ ( .D(n4799), .CLK(CK), .RSTB(n5240), .Q(
        n5008), .QN(n846) );
  DFFARX1_RVT InstQueue_reg_10__1_ ( .D(n4807), .CLK(CK), .RSTB(n5240), .Q(
        n5006), .QN(n854) );
  DFFARX1_RVT InstQueue_reg_9__1_ ( .D(n4815), .CLK(CK), .RSTB(n5240), .Q(
        n5005), .QN(n862) );
  DFFARX1_RVT InstQueue_reg_8__1_ ( .D(n4823), .CLK(CK), .RSTB(n5240), .Q(
        n5140), .QN(n870) );
  DFFARX1_RVT InstQueue_reg_7__1_ ( .D(n4831), .CLK(CK), .RSTB(n5240), .Q(
        n5009), .QN(n878) );
  DFFARX1_RVT InstQueue_reg_6__1_ ( .D(n4839), .CLK(CK), .RSTB(n5240), .Q(
        n5007), .QN(n886) );
  DFFARX1_RVT InstQueue_reg_5__1_ ( .D(n4847), .CLK(CK), .RSTB(n5240), .Q(
        n5004), .QN(n894) );
  DFFARX1_RVT InstQueue_reg_4__1_ ( .D(n4855), .CLK(CK), .RSTB(n5240), .Q(
        n5139), .QN(n902) );
  DFFARX1_RVT InstQueue_reg_3__1_ ( .D(n4863), .CLK(CK), .RSTB(n5239), .Q(
        n5141), .QN(n910) );
  DFFARX1_RVT InstQueue_reg_2__1_ ( .D(n4871), .CLK(CK), .RSTB(n5239), .Q(
        n5137), .QN(n918) );
  DFFARX1_RVT InstQueue_reg_1__1_ ( .D(n4879), .CLK(CK), .RSTB(n5239), .Q(
        n5129), .QN(n926) );
  DFFARX1_RVT InstQueue_reg_0__1_ ( .D(n4887), .CLK(CK), .RSTB(n5246), .Q(
        n5128), .QN(n934) );
  DFFARX1_RVT InstQueue_reg_15__0_ ( .D(n4768), .CLK(CK), .RSTB(n5236), .QN(
        n815) );
  DFFARX1_RVT InstQueue_reg_14__0_ ( .D(n4776), .CLK(CK), .RSTB(n5236), .Q(
        n5117), .QN(n823) );
  DFFARX1_RVT InstQueue_reg_13__0_ ( .D(n4784), .CLK(CK), .RSTB(n5236), .Q(
        n4996), .QN(n831) );
  DFFARX1_RVT InstQueue_reg_12__0_ ( .D(n4792), .CLK(CK), .RSTB(n5236), .Q(
        n5133), .QN(n839) );
  DFFARX1_RVT InstQueue_reg_11__0_ ( .D(n4800), .CLK(CK), .RSTB(n5236), .Q(
        n5001), .QN(n847) );
  DFFARX1_RVT InstQueue_reg_10__0_ ( .D(n4808), .CLK(CK), .RSTB(n5247), .Q(
        n4999), .QN(n855) );
  DFFARX1_RVT InstQueue_reg_9__0_ ( .D(n4816), .CLK(CK), .RSTB(n5236), .Q(
        n4998), .QN(n863) );
  DFFARX1_RVT InstQueue_reg_8__0_ ( .D(n4824), .CLK(CK), .RSTB(n5236), .Q(
        n5135), .QN(n871) );
  DFFARX1_RVT InstQueue_reg_7__0_ ( .D(n4832), .CLK(CK), .RSTB(n5236), .Q(
        n5002), .QN(n879) );
  DFFARX1_RVT InstQueue_reg_6__0_ ( .D(n4840), .CLK(CK), .RSTB(n5236), .Q(
        n5000), .QN(n887) );
  DFFARX1_RVT InstQueue_reg_5__0_ ( .D(n4848), .CLK(CK), .RSTB(n5235), .Q(
        n4997), .QN(n895) );
  DFFARX1_RVT InstQueue_reg_4__0_ ( .D(n4856), .CLK(CK), .RSTB(n5235), .Q(
        n5134), .QN(n903) );
  DFFARX1_RVT InstQueue_reg_3__0_ ( .D(n4864), .CLK(CK), .RSTB(n5235), .Q(
        n5136), .QN(n911) );
  DFFARX1_RVT InstQueue_reg_2__0_ ( .D(n4872), .CLK(CK), .RSTB(n5235), .Q(
        n5132), .QN(n919) );
  DFFARX1_RVT InstQueue_reg_1__0_ ( .D(n4880), .CLK(CK), .RSTB(n5235), .Q(
        n5123), .QN(n927) );
  DFFARX1_RVT InstQueue_reg_0__0_ ( .D(n4888), .CLK(CK), .RSTB(n5235), .Q(
        n5118), .QN(n935) );
  DFFARX1_RVT InstQueue_reg_0__4_ ( .D(n4884), .CLK(CK), .RSTB(n5246), .Q(
        n5120), .QN(n931) );
  DFFARX1_RVT InstQueue_reg_1__4_ ( .D(n4876), .CLK(CK), .RSTB(n5241), .Q(
        n5125), .QN(n923) );
  DFFARX1_RVT InstQueue_reg_2__4_ ( .D(n4868), .CLK(CK), .RSTB(n5241), .Q(
        n5152), .QN(n915) );
  DFFARX1_RVT InstQueue_reg_3__4_ ( .D(n4860), .CLK(CK), .RSTB(n5241), .Q(
        n5156), .QN(n907) );
  DFFARX1_RVT InstQueue_reg_4__4_ ( .D(n4852), .CLK(CK), .RSTB(n5241), .Q(
        n5154), .QN(n899) );
  DFFARX1_RVT InstQueue_reg_5__4_ ( .D(n4844), .CLK(CK), .RSTB(n5241), .Q(
        n5024), .QN(n891) );
  DFFARX1_RVT InstQueue_reg_6__4_ ( .D(n4836), .CLK(CK), .RSTB(n5241), .Q(
        n5027), .QN(n883) );
  DFFARX1_RVT InstQueue_reg_7__4_ ( .D(n4828), .CLK(CK), .RSTB(n5241), .Q(
        n5029), .QN(n875) );
  DFFARX1_RVT InstQueue_reg_8__4_ ( .D(n4820), .CLK(CK), .RSTB(n5241), .Q(
        n5155), .QN(n867) );
  DFFARX1_RVT InstQueue_reg_9__4_ ( .D(n4812), .CLK(CK), .RSTB(n5241), .Q(
        n5025), .QN(n859) );
  DFFARX1_RVT InstQueue_reg_10__4_ ( .D(n4804), .CLK(CK), .RSTB(n5241), .Q(
        n5026), .QN(n851) );
  DFFARX1_RVT InstQueue_reg_11__4_ ( .D(n4796), .CLK(CK), .RSTB(n5241), .Q(
        n5028), .QN(n843) );
  DFFARX1_RVT InstQueue_reg_12__4_ ( .D(n4788), .CLK(CK), .RSTB(n5241), .Q(
        n5153), .QN(n835) );
  DFFARX1_RVT InstQueue_reg_13__4_ ( .D(n4780), .CLK(CK), .RSTB(n5242), .Q(
        n5023), .QN(n827) );
  DFFARX1_RVT InstQueue_reg_14__4_ ( .D(n4772), .CLK(CK), .RSTB(n5242), .Q(
        n5115), .QN(n819) );
  DFFARX1_RVT InstQueue_reg_15__4_ ( .D(n4764), .CLK(CK), .RSTB(n5242), .QN(
        n807) );
  DFFARX1_RVT InstQueue_reg_15__5_ ( .D(n4763), .CLK(CK), .RSTB(n5243), .QN(
        n805) );
  DFFARX1_RVT InstQueue_reg_14__5_ ( .D(n4771), .CLK(CK), .RSTB(n5243), .Q(
        n5116), .QN(n818) );
  DFFARX1_RVT InstQueue_reg_13__5_ ( .D(n4779), .CLK(CK), .RSTB(n5243), .Q(
        n5030), .QN(n826) );
  DFFARX1_RVT InstQueue_reg_12__5_ ( .D(n4787), .CLK(CK), .RSTB(n5243), .Q(
        n5158), .QN(n834) );
  DFFARX1_RVT InstQueue_reg_11__5_ ( .D(n4795), .CLK(CK), .RSTB(n5243), .Q(
        n5035), .QN(n842) );
  DFFARX1_RVT InstQueue_reg_10__5_ ( .D(n4803), .CLK(CK), .RSTB(n5243), .Q(
        n5033), .QN(n850) );
  DFFARX1_RVT InstQueue_reg_9__5_ ( .D(n4811), .CLK(CK), .RSTB(n5242), .Q(
        n5032), .QN(n858) );
  DFFARX1_RVT InstQueue_reg_8__5_ ( .D(n4819), .CLK(CK), .RSTB(n5242), .Q(
        n5160), .QN(n866) );
  DFFARX1_RVT InstQueue_reg_7__5_ ( .D(n4827), .CLK(CK), .RSTB(n5242), .Q(
        n5036), .QN(n874) );
  DFFARX1_RVT InstQueue_reg_6__5_ ( .D(n4835), .CLK(CK), .RSTB(n5242), .Q(
        n5034), .QN(n882) );
  DFFARX1_RVT InstQueue_reg_5__5_ ( .D(n4843), .CLK(CK), .RSTB(n5242), .Q(
        n5031), .QN(n890) );
  DFFARX1_RVT InstQueue_reg_4__5_ ( .D(n4851), .CLK(CK), .RSTB(n5242), .Q(
        n5159), .QN(n898) );
  DFFARX1_RVT InstQueue_reg_3__5_ ( .D(n4859), .CLK(CK), .RSTB(n5242), .Q(
        n5161), .QN(n906) );
  DFFARX1_RVT InstQueue_reg_2__5_ ( .D(n4867), .CLK(CK), .RSTB(n5242), .Q(
        n5157), .QN(n914) );
  DFFARX1_RVT InstQueue_reg_1__5_ ( .D(n4875), .CLK(CK), .RSTB(n5242), .Q(
        n5126), .QN(n922) );
  DFFARX1_RVT InstQueue_reg_0__5_ ( .D(n4883), .CLK(CK), .RSTB(n5243), .Q(
        n5121), .QN(n930) );
  DFFARX1_RVT InstQueue_reg_15__6_ ( .D(n4762), .CLK(CK), .RSTB(n5246), .QN(
        n803) );
  DFFARX1_RVT InstQueue_reg_14__6_ ( .D(n4770), .CLK(CK), .RSTB(n5246), .Q(
        n5111), .QN(n817) );
  DFFARX1_RVT InstQueue_reg_13__6_ ( .D(n4778), .CLK(CK), .RSTB(n5245), .Q(
        n5037), .QN(n825) );
  DFFARX1_RVT InstQueue_reg_12__6_ ( .D(n4786), .CLK(CK), .RSTB(n5245), .Q(
        n5163), .QN(n833) );
  DFFARX1_RVT InstQueue_reg_11__6_ ( .D(n4794), .CLK(CK), .RSTB(n5245), .Q(
        n5042), .QN(n841) );
  DFFARX1_RVT InstQueue_reg_10__6_ ( .D(n4802), .CLK(CK), .RSTB(n5245), .Q(
        n5040), .QN(n849) );
  DFFARX1_RVT InstQueue_reg_9__6_ ( .D(n4810), .CLK(CK), .RSTB(n5245), .Q(
        n5039), .QN(n857) );
  DFFARX1_RVT InstQueue_reg_8__6_ ( .D(n4818), .CLK(CK), .RSTB(n5245), .Q(
        n5165), .QN(n865) );
  DFFARX1_RVT InstQueue_reg_7__6_ ( .D(n4826), .CLK(CK), .RSTB(n5245), .Q(
        n5109), .QN(n873) );
  DFFARX1_RVT InstQueue_reg_6__6_ ( .D(n4834), .CLK(CK), .RSTB(n5245), .Q(
        n5041), .QN(n881) );
  DFFARX1_RVT InstQueue_reg_5__6_ ( .D(n4842), .CLK(CK), .RSTB(n5245), .Q(
        n5038), .QN(n889) );
  DFFARX1_RVT InstQueue_reg_4__6_ ( .D(n4850), .CLK(CK), .RSTB(n5245), .Q(
        n5164), .QN(n897) );
  DFFARX1_RVT InstQueue_reg_3__6_ ( .D(n4858), .CLK(CK), .RSTB(n5245), .Q(
        n5166), .QN(n905) );
  DFFARX1_RVT InstQueue_reg_2__6_ ( .D(n4866), .CLK(CK), .RSTB(n5245), .Q(
        n5162), .QN(n913) );
  DFFARX1_RVT InstQueue_reg_1__6_ ( .D(n4874), .CLK(CK), .RSTB(n5244), .Q(
        n5127), .QN(n921) );
  DFFARX1_RVT InstQueue_reg_0__6_ ( .D(n4882), .CLK(CK), .RSTB(n5246), .Q(
        n5122), .QN(n929) );
  DFFARX1_RVT ReadRequest_reg ( .D(n4721), .CLK(CK), .RSTB(n5239), .QN(n9512)
         );
  DFFARX1_RVT W_R_n_reg ( .D(n4720), .CLK(CK), .RSTB(n5239), .Q(W_R_n) );
  DFFARX1_RVT More_reg ( .D(n4722), .CLK(CK), .RSTB(n5219), .QN(n9513) );
  DFFARX1_RVT EBX_reg_30_ ( .D(n4622), .CLK(CK), .RSTB(n5220), .Q(n4988), .QN(
        n9521) );
  DFFARX1_RVT EBX_reg_29_ ( .D(n4623), .CLK(CK), .RSTB(n5220), .Q(n4980), .QN(
        n9523) );
  DFFARX1_RVT EBX_reg_28_ ( .D(n4624), .CLK(CK), .RSTB(n5220), .Q(n4981), .QN(
        n9524) );
  DFFARX1_RVT EBX_reg_27_ ( .D(n4625), .CLK(CK), .RSTB(n5221), .Q(n4982), .QN(
        n9525) );
  DFFARX1_RVT EBX_reg_26_ ( .D(n4626), .CLK(CK), .RSTB(n5221), .Q(n4983), .QN(
        n9526) );
  DFFARX1_RVT EBX_reg_25_ ( .D(n4627), .CLK(CK), .RSTB(n5221), .Q(n4984), .QN(
        n9527) );
  DFFARX1_RVT EBX_reg_24_ ( .D(n4628), .CLK(CK), .RSTB(n5222), .Q(n4985), .QN(
        n9528) );
  DFFARX1_RVT EBX_reg_23_ ( .D(n4629), .CLK(CK), .RSTB(n5222), .Q(n4990), .QN(
        n9529) );
  DFFARX1_RVT EBX_reg_22_ ( .D(n4630), .CLK(CK), .RSTB(n5222), .Q(n4991), .QN(
        n9530) );
  DFFARX1_RVT EBX_reg_21_ ( .D(n4631), .CLK(CK), .RSTB(n5223), .Q(n4995), .QN(
        n9531) );
  DFFARX1_RVT EBX_reg_20_ ( .D(n4632), .CLK(CK), .RSTB(n5223), .Q(n4994), .QN(
        n9532) );
  DFFARX1_RVT EBX_reg_19_ ( .D(n4633), .CLK(CK), .RSTB(n5223), .Q(n4993), .QN(
        n9534) );
  DFFARX1_RVT EBX_reg_18_ ( .D(n4634), .CLK(CK), .RSTB(n5224), .Q(n4992), .QN(
        n9535) );
  DFFARX1_RVT EBX_reg_17_ ( .D(n4635), .CLK(CK), .RSTB(n5224), .Q(n4987), .QN(
        n9536) );
  DFFARX1_RVT EBX_reg_16_ ( .D(n4636), .CLK(CK), .RSTB(n5224), .Q(n4986), .QN(
        n9537) );
  DFFARX1_RVT EBX_reg_15_ ( .D(n4637), .CLK(CK), .RSTB(n5225), .Q(n4932), .QN(
        n9538) );
  DFFARX1_RVT EBX_reg_14_ ( .D(n4638), .CLK(CK), .RSTB(n5225), .Q(n4934), .QN(
        n9539) );
  DFFARX1_RVT EBX_reg_13_ ( .D(n4639), .CLK(CK), .RSTB(n5227), .Q(n4935), .QN(
        n9540) );
  DFFARX1_RVT EBX_reg_12_ ( .D(n4640), .CLK(CK), .RSTB(n5227), .Q(n4944), .QN(
        n9541) );
  DFFARX1_RVT EBX_reg_11_ ( .D(n4641), .CLK(CK), .RSTB(n5227), .Q(n4936), .QN(
        n9542) );
  DFFARX1_RVT EBX_reg_10_ ( .D(n4642), .CLK(CK), .RSTB(n5228), .Q(n4966) );
  DFFARX1_RVT EBX_reg_9_ ( .D(n4643), .CLK(CK), .RSTB(n5228), .Q(n4933), .QN(
        n9515) );
  DFFARX1_RVT EBX_reg_8_ ( .D(n4644), .CLK(CK), .RSTB(n5228), .Q(n4943), .QN(
        n9516) );
  DFFARX1_RVT EBX_reg_7_ ( .D(n4645), .CLK(CK), .RSTB(n5229), .Q(n4937), .QN(
        n9517) );
  DFFARX1_RVT EBX_reg_6_ ( .D(n4646), .CLK(CK), .RSTB(n5229), .Q(n4942), .QN(
        n9518) );
  DFFARX1_RVT EBX_reg_5_ ( .D(n4647), .CLK(CK), .RSTB(n5229), .Q(n4938), .QN(
        n9519) );
  DFFARX1_RVT EBX_reg_4_ ( .D(n4648), .CLK(CK), .RSTB(n5230), .Q(n4941), .QN(
        n9520) );
  DFFARX1_RVT EBX_reg_3_ ( .D(n4649), .CLK(CK), .RSTB(n5230), .Q(n4939), .QN(
        n9522) );
  DFFARX1_RVT EBX_reg_2_ ( .D(n4650), .CLK(CK), .RSTB(n5231), .Q(n4940), .QN(
        n9533) );
  DFFARX1_RVT EBX_reg_1_ ( .D(n4651), .CLK(CK), .RSTB(n5231), .Q(n4964), .QN(
        n9543) );
  DFFARX1_RVT EBX_reg_0_ ( .D(n4652), .CLK(CK), .RSTB(n5235), .Q(n4911), .QN(
        n9544) );
  DFFARX1_RVT InstQueue_reg_15__7_ ( .D(n4894), .CLK(CK), .RSTB(n5244), .Q(
        n5194), .QN(n801) );
  DFFARX1_RVT InstQueue_reg_0__7_ ( .D(n4881), .CLK(CK), .RSTB(n5243), .Q(
        n5049), .QN(n928) );
  DFFARX1_RVT InstQueue_reg_1__7_ ( .D(n4873), .CLK(CK), .RSTB(n5243), .Q(
        n5167), .QN(n920) );
  DFFARX1_RVT InstQueue_reg_2__7_ ( .D(n4865), .CLK(CK), .RSTB(n5243), .Q(
        n5168), .QN(n912) );
  DFFARX1_RVT InstQueue_reg_3__7_ ( .D(n4857), .CLK(CK), .RSTB(n5243), .Q(
        n5172), .QN(n904) );
  DFFARX1_RVT InstQueue_reg_4__7_ ( .D(n4849), .CLK(CK), .RSTB(n5243), .Q(
        n5169), .QN(n896) );
  DFFARX1_RVT InstQueue_reg_5__7_ ( .D(n4841), .CLK(CK), .RSTB(n5244), .Q(
        n5043), .QN(n888) );
  DFFARX1_RVT InstQueue_reg_6__7_ ( .D(n4833), .CLK(CK), .RSTB(n5244), .Q(
        n5046), .QN(n880) );
  DFFARX1_RVT InstQueue_reg_7__7_ ( .D(n4825), .CLK(CK), .RSTB(n5244), .Q(
        n5050), .QN(n872) );
  DFFARX1_RVT InstQueue_reg_8__7_ ( .D(n4817), .CLK(CK), .RSTB(n5244), .Q(
        n5170), .QN(n864) );
  DFFARX1_RVT InstQueue_reg_9__7_ ( .D(n4809), .CLK(CK), .RSTB(n5244), .Q(
        n5044), .QN(n856) );
  DFFARX1_RVT InstQueue_reg_10__7_ ( .D(n4801), .CLK(CK), .RSTB(n5244), .Q(
        n5047), .QN(n848) );
  DFFARX1_RVT InstQueue_reg_11__7_ ( .D(n4793), .CLK(CK), .RSTB(n5244), .Q(
        n5051), .QN(n840) );
  DFFARX1_RVT InstQueue_reg_12__7_ ( .D(n4785), .CLK(CK), .RSTB(n5244), .Q(
        n5171), .QN(n832) );
  DFFARX1_RVT InstQueue_reg_13__7_ ( .D(n4777), .CLK(CK), .RSTB(n5244), .Q(
        n5045), .QN(n824) );
  DFFARX1_RVT lWord_reg_0_ ( .D(n4699), .CLK(CK), .RSTB(n5235), .Q(n5176) );
  DFFARX1_RVT EAX_reg_0_ ( .D(n4715), .CLK(CK), .RSTB(n5235), .Q(n4961), .QN(
        n9560) );
  DFFARX1_RVT uWord_reg_0_ ( .D(n4667), .CLK(CK), .RSTB(n5235), .Q(uWord[0])
         );
  DFFARX1_RVT Datao_reg_0_ ( .D(n4526), .CLK(CK), .RSTB(n5235), .Q(Datao[0])
         );
  DFFARX1_RVT EAX_reg_1_ ( .D(n4714), .CLK(CK), .RSTB(n5231), .Q(n4959), .QN(
        n9559) );
  DFFARX1_RVT lWord_reg_1_ ( .D(n4698), .CLK(CK), .RSTB(n5226), .Q(n5175) );
  DFFARX1_RVT uWord_reg_1_ ( .D(n4666), .CLK(CK), .RSTB(n5231), .Q(uWord[1])
         );
  DFFARX1_RVT Datao_reg_1_ ( .D(n4525), .CLK(CK), .RSTB(n5226), .Q(Datao[1])
         );
  DFFARX1_RVT EAX_reg_2_ ( .D(n4713), .CLK(CK), .RSTB(n5234), .Q(n4957), .QN(
        n9552) );
  DFFARX1_RVT lWord_reg_2_ ( .D(n4697), .CLK(CK), .RSTB(n5234), .Q(n5177) );
  DFFARX1_RVT uWord_reg_2_ ( .D(n4665), .CLK(CK), .RSTB(n5234), .Q(uWord[2])
         );
  DFFARX1_RVT Datao_reg_2_ ( .D(n4524), .CLK(CK), .RSTB(n5231), .Q(Datao[2])
         );
  DFFARX1_RVT EAX_reg_3_ ( .D(n4712), .CLK(CK), .RSTB(n5234), .Q(n4951), .QN(
        n9551) );
  DFFARX1_RVT lWord_reg_3_ ( .D(n4696), .CLK(CK), .RSTB(n5234), .Q(n5178) );
  DFFARX1_RVT uWord_reg_3_ ( .D(n4664), .CLK(CK), .RSTB(n5234), .Q(uWord[3])
         );
  DFFARX1_RVT Datao_reg_3_ ( .D(n4523), .CLK(CK), .RSTB(n5230), .Q(Datao[3])
         );
  DFFARX1_RVT EAX_reg_4_ ( .D(n4711), .CLK(CK), .RSTB(n5234), .Q(n4954), .QN(
        n9550) );
  DFFARX1_RVT lWord_reg_4_ ( .D(n4695), .CLK(CK), .RSTB(n5234), .Q(n5179) );
  DFFARX1_RVT uWord_reg_4_ ( .D(n4663), .CLK(CK), .RSTB(n5234), .Q(uWord[4])
         );
  DFFARX1_RVT Datao_reg_4_ ( .D(n4522), .CLK(CK), .RSTB(n5230), .Q(Datao[4])
         );
  DFFARX1_RVT EAX_reg_5_ ( .D(n4710), .CLK(CK), .RSTB(n5234), .Q(n4948), .QN(
        n9549) );
  DFFARX1_RVT lWord_reg_5_ ( .D(n4694), .CLK(CK), .RSTB(n5233), .Q(n5180) );
  DFFARX1_RVT uWord_reg_5_ ( .D(n4662), .CLK(CK), .RSTB(n5234), .Q(uWord[5])
         );
  DFFARX1_RVT Datao_reg_5_ ( .D(n4521), .CLK(CK), .RSTB(n5229), .Q(Datao[5])
         );
  DFFARX1_RVT EAX_reg_6_ ( .D(n4709), .CLK(CK), .RSTB(n5233), .Q(n4956), .QN(
        n9548) );
  DFFARX1_RVT lWord_reg_6_ ( .D(n4693), .CLK(CK), .RSTB(n5233), .Q(n5181) );
  DFFARX1_RVT uWord_reg_6_ ( .D(n4661), .CLK(CK), .RSTB(n5233), .Q(uWord[6])
         );
  DFFARX1_RVT Datao_reg_6_ ( .D(n4520), .CLK(CK), .RSTB(n5229), .Q(Datao[6])
         );
  DFFARX1_RVT EAX_reg_7_ ( .D(n4708), .CLK(CK), .RSTB(n5233), .Q(n4950), .QN(
        n9547) );
  DFFARX1_RVT lWord_reg_7_ ( .D(n4692), .CLK(CK), .RSTB(n5233), .Q(n5182) );
  DFFARX1_RVT uWord_reg_7_ ( .D(n4660), .CLK(CK), .RSTB(n5233), .Q(uWord[7])
         );
  DFFARX1_RVT Datao_reg_7_ ( .D(n4519), .CLK(CK), .RSTB(n5229), .Q(Datao[7])
         );
  DFFARX1_RVT EAX_reg_8_ ( .D(n4707), .CLK(CK), .RSTB(n5233), .Q(n4953), .QN(
        n9546) );
  DFFARX1_RVT lWord_reg_8_ ( .D(n4691), .CLK(CK), .RSTB(n5233), .Q(n5183) );
  DFFARX1_RVT uWord_reg_8_ ( .D(n4659), .CLK(CK), .RSTB(n5233), .Q(uWord[8])
         );
  DFFARX1_RVT Datao_reg_8_ ( .D(n4518), .CLK(CK), .RSTB(n5228), .Q(Datao[8])
         );
  DFFARX1_RVT EAX_reg_9_ ( .D(n4706), .CLK(CK), .RSTB(n5233), .Q(n4947), .QN(
        n9545) );
  DFFARX1_RVT lWord_reg_9_ ( .D(n4690), .CLK(CK), .RSTB(n5232), .Q(n5184) );
  DFFARX1_RVT uWord_reg_9_ ( .D(n4658), .CLK(CK), .RSTB(n5233), .Q(uWord[9])
         );
  DFFARX1_RVT Datao_reg_9_ ( .D(n4517), .CLK(CK), .RSTB(n5228), .Q(Datao[9])
         );
  DFFARX1_RVT EAX_reg_10_ ( .D(n4705), .CLK(CK), .RSTB(n5232), .Q(n4952), .QN(
        n9558) );
  DFFARX1_RVT lWord_reg_10_ ( .D(n4689), .CLK(CK), .RSTB(n5232), .Q(n5185) );
  DFFARX1_RVT uWord_reg_10_ ( .D(n4657), .CLK(CK), .RSTB(n5232), .Q(uWord[10])
         );
  DFFARX1_RVT Datao_reg_10_ ( .D(n4516), .CLK(CK), .RSTB(n5228), .Q(Datao[10])
         );
  DFFARX1_RVT EAX_reg_11_ ( .D(n4704), .CLK(CK), .RSTB(n5232), .Q(n4946), .QN(
        n9557) );
  DFFARX1_RVT lWord_reg_11_ ( .D(n4688), .CLK(CK), .RSTB(n5232), .Q(n5186) );
  DFFARX1_RVT uWord_reg_11_ ( .D(n4656), .CLK(CK), .RSTB(n5232), .Q(uWord[11])
         );
  DFFARX1_RVT Datao_reg_11_ ( .D(n4515), .CLK(CK), .RSTB(n5227), .Q(Datao[11])
         );
  DFFARX1_RVT EAX_reg_12_ ( .D(n4703), .CLK(CK), .RSTB(n5232), .Q(n4955), .QN(
        n9556) );
  DFFARX1_RVT lWord_reg_12_ ( .D(n4687), .CLK(CK), .RSTB(n5232), .Q(n5187) );
  DFFARX1_RVT uWord_reg_12_ ( .D(n4655), .CLK(CK), .RSTB(n5232), .Q(uWord[12])
         );
  DFFARX1_RVT Datao_reg_12_ ( .D(n4514), .CLK(CK), .RSTB(n5227), .Q(Datao[12])
         );
  DFFARX1_RVT EAX_reg_13_ ( .D(n4702), .CLK(CK), .RSTB(n5232), .Q(n4949), .QN(
        n9555) );
  DFFARX1_RVT lWord_reg_13_ ( .D(n4686), .CLK(CK), .RSTB(n5231), .Q(n5188) );
  DFFARX1_RVT uWord_reg_13_ ( .D(n4654), .CLK(CK), .RSTB(n5232), .Q(uWord[13])
         );
  DFFARX1_RVT Datao_reg_13_ ( .D(n4513), .CLK(CK), .RSTB(n5227), .Q(Datao[13])
         );
  DFFARX1_RVT EAX_reg_14_ ( .D(n4701), .CLK(CK), .RSTB(n5225), .Q(n4960), .QN(
        n9554) );
  DFFARX1_RVT lWord_reg_14_ ( .D(n4685), .CLK(CK), .RSTB(n5219), .Q(n5189) );
  DFFARX1_RVT uWord_reg_14_ ( .D(n4653), .CLK(CK), .RSTB(n5225), .Q(uWord[14])
         );
  DFFARX1_RVT Datao_reg_14_ ( .D(n4512), .CLK(CK), .RSTB(n5219), .Q(Datao[14])
         );
  DFFARX1_RVT EAX_reg_15_ ( .D(n4700), .CLK(CK), .RSTB(n5231), .Q(n4945), .QN(
        n9553) );
  DFFARX1_RVT lWord_reg_15_ ( .D(n4684), .CLK(CK), .RSTB(n5219), .Q(n5174) );
  DFFARX1_RVT Datao_reg_15_ ( .D(n4511), .CLK(CK), .RSTB(n5219), .Q(Datao[15])
         );
  DFFARX1_RVT EAX_reg_16_ ( .D(n4683), .CLK(CK), .RSTB(n5234), .Q(n5088) );
  DFFARX1_RVT Datao_reg_16_ ( .D(n4510), .CLK(CK), .RSTB(n5224), .Q(Datao[16])
         );
  DFFARX1_RVT EAX_reg_17_ ( .D(n4682), .CLK(CK), .RSTB(n5231), .Q(n5087) );
  DFFARX1_RVT Datao_reg_17_ ( .D(n4509), .CLK(CK), .RSTB(n5224), .Q(Datao[17])
         );
  DFFARX1_RVT EAX_reg_18_ ( .D(n4681), .CLK(CK), .RSTB(n5226), .Q(n5089) );
  DFFARX1_RVT Datao_reg_18_ ( .D(n4508), .CLK(CK), .RSTB(n5224), .Q(Datao[18])
         );
  DFFARX1_RVT EAX_reg_19_ ( .D(n4680), .CLK(CK), .RSTB(n5226), .Q(n5090) );
  DFFARX1_RVT Datao_reg_19_ ( .D(n4507), .CLK(CK), .RSTB(n5223), .Q(Datao[19])
         );
  DFFARX1_RVT EAX_reg_20_ ( .D(n4679), .CLK(CK), .RSTB(n5226), .Q(n5091) );
  DFFARX1_RVT Datao_reg_20_ ( .D(n4506), .CLK(CK), .RSTB(n5223), .Q(Datao[20])
         );
  DFFARX1_RVT EAX_reg_21_ ( .D(n4678), .CLK(CK), .RSTB(n5226), .Q(n5092) );
  DFFARX1_RVT Datao_reg_21_ ( .D(n4505), .CLK(CK), .RSTB(n5223), .Q(Datao[21])
         );
  DFFARX1_RVT EAX_reg_22_ ( .D(n4677), .CLK(CK), .RSTB(n5226), .Q(n5093) );
  DFFARX1_RVT Datao_reg_22_ ( .D(n4504), .CLK(CK), .RSTB(n5222), .Q(Datao[22])
         );
  DFFARX1_RVT EAX_reg_23_ ( .D(n4676), .CLK(CK), .RSTB(n5226), .Q(n5094) );
  DFFARX1_RVT Datao_reg_23_ ( .D(n4503), .CLK(CK), .RSTB(n5222), .Q(Datao[23])
         );
  DFFARX1_RVT EAX_reg_24_ ( .D(n4675), .CLK(CK), .RSTB(n5226), .Q(n5095) );
  DFFARX1_RVT Datao_reg_24_ ( .D(n4502), .CLK(CK), .RSTB(n5222), .Q(Datao[24])
         );
  DFFARX1_RVT EAX_reg_25_ ( .D(n4674), .CLK(CK), .RSTB(n5226), .Q(n5096) );
  DFFARX1_RVT Datao_reg_25_ ( .D(n4501), .CLK(CK), .RSTB(n5221), .Q(Datao[25])
         );
  DFFARX1_RVT EAX_reg_26_ ( .D(n4673), .CLK(CK), .RSTB(n5225), .Q(n5097) );
  DFFARX1_RVT Datao_reg_26_ ( .D(n4500), .CLK(CK), .RSTB(n5221), .Q(Datao[26])
         );
  DFFARX1_RVT EAX_reg_27_ ( .D(n4672), .CLK(CK), .RSTB(n5225), .Q(n5098) );
  DFFARX1_RVT Datao_reg_27_ ( .D(n4499), .CLK(CK), .RSTB(n5221), .Q(Datao[27])
         );
  DFFARX1_RVT EAX_reg_28_ ( .D(n4671), .CLK(CK), .RSTB(n5225), .Q(n5099) );
  DFFARX1_RVT Datao_reg_28_ ( .D(n4498), .CLK(CK), .RSTB(n5220), .Q(Datao[28])
         );
  DFFARX1_RVT EAX_reg_29_ ( .D(n4670), .CLK(CK), .RSTB(n5225), .Q(n5100) );
  DFFARX1_RVT Datao_reg_29_ ( .D(n4497), .CLK(CK), .RSTB(n5220), .Q(Datao[29])
         );
  DFFARX1_RVT EAX_reg_30_ ( .D(n4669), .CLK(CK), .RSTB(n5225), .Q(n5101) );
  DFFARX1_RVT EAX_reg_31_ ( .D(n4668), .CLK(CK), .RSTB(n5219), .Q(n5054) );
  DFFARX1_RVT PhyAddrPointer_reg_1_ ( .D(n4557), .CLK(CK), .RSTB(n5231), .Q(
        n5063) );
  DFFARX1_RVT rEIP_reg_1_ ( .D(n4619), .CLK(CK), .RSTB(n5231), .Q(rEIP[1]), 
        .QN(n5053) );
  DFFARX1_RVT InstAddrPointer_reg_1_ ( .D(n4723), .CLK(CK), .RSTB(n5231), .Q(
        n5052), .QN(n9575) );
  DFFARX1_RVT PhyAddrPointer_reg_2_ ( .D(n4556), .CLK(CK), .RSTB(n5230), .Q(
        n5062) );
  DFFARX1_RVT rEIP_reg_2_ ( .D(n4618), .CLK(CK), .RSTB(n5231), .Q(rEIP[2]) );
  DFFARX1_RVT InstAddrPointer_reg_2_ ( .D(n4724), .CLK(CK), .RSTB(n5230), .Q(
        n5107), .QN(n9569) );
  DFFARX1_RVT PhyAddrPointer_reg_3_ ( .D(n4555), .CLK(CK), .RSTB(n5230), .Q(
        n5061) );
  DFFARX1_RVT rEIP_reg_3_ ( .D(n4617), .CLK(CK), .RSTB(n5230), .Q(rEIP[3]) );
  DFFARX1_RVT InstAddrPointer_reg_3_ ( .D(n4725), .CLK(CK), .RSTB(n5230), .Q(
        n5106), .QN(n9566) );
  DFFARX1_RVT PhyAddrPointer_reg_4_ ( .D(n4554), .CLK(CK), .RSTB(n5230), .Q(
        n5060) );
  DFFARX1_RVT rEIP_reg_4_ ( .D(n4616), .CLK(CK), .RSTB(n5230), .Q(rEIP[4]) );
  DFFARX1_RVT InstAddrPointer_reg_4_ ( .D(n4726), .CLK(CK), .RSTB(n5230), .Q(
        n5105), .QN(n9565) );
  DFFARX1_RVT PhyAddrPointer_reg_5_ ( .D(n4553), .CLK(CK), .RSTB(n5229), .Q(
        n5059) );
  DFFARX1_RVT rEIP_reg_5_ ( .D(n4615), .CLK(CK), .RSTB(n5229), .Q(rEIP[5]) );
  DFFARX1_RVT InstAddrPointer_reg_5_ ( .D(n4727), .CLK(CK), .RSTB(n5229), .Q(
        n5104), .QN(n9564) );
  DFFARX1_RVT PhyAddrPointer_reg_6_ ( .D(n4552), .CLK(CK), .RSTB(n5229), .Q(
        n5058) );
  DFFARX1_RVT rEIP_reg_6_ ( .D(n4614), .CLK(CK), .RSTB(n5229), .Q(rEIP[6]) );
  DFFARX1_RVT InstAddrPointer_reg_6_ ( .D(n4728), .CLK(CK), .RSTB(n5229), .Q(
        n5103), .QN(n9563) );
  DFFARX1_RVT PhyAddrPointer_reg_7_ ( .D(n4551), .CLK(CK), .RSTB(n5228), .Q(
        n5057) );
  DFFARX1_RVT rEIP_reg_7_ ( .D(n4613), .CLK(CK), .RSTB(n5228), .Q(rEIP[7]) );
  DFFARX1_RVT InstAddrPointer_reg_7_ ( .D(n4729), .CLK(CK), .RSTB(n5249), .Q(
        n5102), .QN(n9562) );
  DFFARX1_RVT PhyAddrPointer_reg_8_ ( .D(n4550), .CLK(CK), .RSTB(n5228), .Q(
        n5064) );
  DFFARX1_RVT rEIP_reg_8_ ( .D(n4612), .CLK(CK), .RSTB(n5228), .Q(rEIP[8]) );
  DFFARX1_RVT InstAddrPointer_reg_8_ ( .D(n4730), .CLK(CK), .RSTB(n5249), .Q(
        n4912) );
  DFFARX1_RVT PhyAddrPointer_reg_9_ ( .D(n4549), .CLK(CK), .RSTB(n5228), .Q(
        n5065) );
  DFFARX1_RVT rEIP_reg_9_ ( .D(n4611), .CLK(CK), .RSTB(n5228), .Q(rEIP[9]) );
  DFFARX1_RVT InstAddrPointer_reg_9_ ( .D(n4731), .CLK(CK), .RSTB(n5249), .Q(
        n4965) );
  DFFARX1_RVT PhyAddrPointer_reg_10_ ( .D(n4548), .CLK(CK), .RSTB(n5227), .Q(
        n5066) );
  DFFARX1_RVT rEIP_reg_10_ ( .D(n4610), .CLK(CK), .RSTB(n5227), .Q(rEIP[10])
         );
  DFFARX1_RVT InstAddrPointer_reg_10_ ( .D(n4732), .CLK(CK), .RSTB(n5249), .Q(
        n4978), .QN(n9580) );
  DFFARX1_RVT PhyAddrPointer_reg_11_ ( .D(n4547), .CLK(CK), .RSTB(n5227), .Q(
        n5067) );
  DFFARX1_RVT rEIP_reg_11_ ( .D(n4609), .CLK(CK), .RSTB(n5227), .Q(rEIP[11])
         );
  DFFARX1_RVT InstAddrPointer_reg_11_ ( .D(n4733), .CLK(CK), .RSTB(n5249), .Q(
        n4924) );
  DFFARX1_RVT PhyAddrPointer_reg_12_ ( .D(n4546), .CLK(CK), .RSTB(n5227), .Q(
        n5068) );
  DFFARX1_RVT rEIP_reg_12_ ( .D(n4608), .CLK(CK), .RSTB(n5227), .Q(rEIP[12])
         );
  DFFARX1_RVT InstAddrPointer_reg_12_ ( .D(n4734), .CLK(CK), .RSTB(n5249), .Q(
        n4977), .QN(n9579) );
  DFFARX1_RVT PhyAddrPointer_reg_13_ ( .D(n4545), .CLK(CK), .RSTB(n5226), .Q(
        n5069) );
  DFFARX1_RVT rEIP_reg_13_ ( .D(n4607), .CLK(CK), .RSTB(n5226), .Q(rEIP[13])
         );
  DFFARX1_RVT InstAddrPointer_reg_13_ ( .D(n4735), .CLK(CK), .RSTB(n5249), .Q(
        n4923) );
  DFFARX1_RVT PhyAddrPointer_reg_14_ ( .D(n4544), .CLK(CK), .RSTB(n5225), .Q(
        n5070) );
  DFFARX1_RVT rEIP_reg_14_ ( .D(n4606), .CLK(CK), .RSTB(n5225), .Q(rEIP[14])
         );
  DFFARX1_RVT InstAddrPointer_reg_14_ ( .D(n4736), .CLK(CK), .RSTB(n5249), .Q(
        n4976), .QN(n9578) );
  DFFARX1_RVT PhyAddrPointer_reg_15_ ( .D(n4543), .CLK(CK), .RSTB(n5224), .Q(
        n5071) );
  DFFARX1_RVT rEIP_reg_15_ ( .D(n4605), .CLK(CK), .RSTB(n5225), .Q(rEIP[15])
         );
  DFFARX1_RVT InstAddrPointer_reg_15_ ( .D(n4737), .CLK(CK), .RSTB(n5248), .Q(
        n4922) );
  DFFARX1_RVT PhyAddrPointer_reg_16_ ( .D(n4542), .CLK(CK), .RSTB(n5224), .Q(
        n5072) );
  DFFARX1_RVT rEIP_reg_16_ ( .D(n4604), .CLK(CK), .RSTB(n5224), .Q(rEIP[16])
         );
  DFFARX1_RVT InstAddrPointer_reg_16_ ( .D(n4738), .CLK(CK), .RSTB(n5248), .Q(
        n4975), .QN(n9577) );
  DFFARX1_RVT PhyAddrPointer_reg_17_ ( .D(n4541), .CLK(CK), .RSTB(n5224), .Q(
        n5073) );
  DFFARX1_RVT rEIP_reg_17_ ( .D(n4603), .CLK(CK), .RSTB(n5224), .Q(rEIP[17])
         );
  DFFARX1_RVT InstAddrPointer_reg_17_ ( .D(n4739), .CLK(CK), .RSTB(n5248), .Q(
        n4921) );
  DFFARX1_RVT PhyAddrPointer_reg_18_ ( .D(n4540), .CLK(CK), .RSTB(n5223), .Q(
        n5074) );
  DFFARX1_RVT rEIP_reg_18_ ( .D(n4602), .CLK(CK), .RSTB(n5224), .Q(rEIP[18])
         );
  DFFARX1_RVT InstAddrPointer_reg_18_ ( .D(n4740), .CLK(CK), .RSTB(n5248), .Q(
        n4974), .QN(n9576) );
  DFFARX1_RVT PhyAddrPointer_reg_19_ ( .D(n4539), .CLK(CK), .RSTB(n5223), .Q(
        n5075) );
  DFFARX1_RVT rEIP_reg_19_ ( .D(n4601), .CLK(CK), .RSTB(n5223), .Q(rEIP[19])
         );
  DFFARX1_RVT InstAddrPointer_reg_19_ ( .D(n4741), .CLK(CK), .RSTB(n5248), .Q(
        n4920) );
  DFFARX1_RVT PhyAddrPointer_reg_20_ ( .D(n4538), .CLK(CK), .RSTB(n5223), .Q(
        n5076) );
  DFFARX1_RVT rEIP_reg_20_ ( .D(n4600), .CLK(CK), .RSTB(n5223), .Q(rEIP[20])
         );
  DFFARX1_RVT InstAddrPointer_reg_20_ ( .D(n4742), .CLK(CK), .RSTB(n5248), .Q(
        n4973), .QN(n9574) );
  DFFARX1_RVT PhyAddrPointer_reg_21_ ( .D(n4537), .CLK(CK), .RSTB(n5222), .Q(
        n5077) );
  DFFARX1_RVT rEIP_reg_21_ ( .D(n4599), .CLK(CK), .RSTB(n5223), .Q(rEIP[21])
         );
  DFFARX1_RVT InstAddrPointer_reg_21_ ( .D(n4743), .CLK(CK), .RSTB(n5248), .Q(
        n4919) );
  DFFARX1_RVT PhyAddrPointer_reg_22_ ( .D(n4536), .CLK(CK), .RSTB(n5222), .Q(
        n5078) );
  DFFARX1_RVT rEIP_reg_22_ ( .D(n4598), .CLK(CK), .RSTB(n5222), .Q(rEIP[22])
         );
  DFFARX1_RVT InstAddrPointer_reg_22_ ( .D(n4744), .CLK(CK), .RSTB(n5248), .Q(
        n4972), .QN(n9573) );
  DFFARX1_RVT PhyAddrPointer_reg_23_ ( .D(n4535), .CLK(CK), .RSTB(n5222), .Q(
        n5079) );
  DFFARX1_RVT rEIP_reg_23_ ( .D(n4597), .CLK(CK), .RSTB(n5222), .Q(rEIP[23])
         );
  DFFARX1_RVT InstAddrPointer_reg_23_ ( .D(n4745), .CLK(CK), .RSTB(n5248), .Q(
        n4918) );
  DFFARX1_RVT PhyAddrPointer_reg_24_ ( .D(n4534), .CLK(CK), .RSTB(n5221), .Q(
        n5080) );
  DFFARX1_RVT rEIP_reg_24_ ( .D(n4596), .CLK(CK), .RSTB(n5222), .Q(rEIP[24])
         );
  DFFARX1_RVT InstAddrPointer_reg_24_ ( .D(n4746), .CLK(CK), .RSTB(n5248), .Q(
        n4971), .QN(n9572) );
  DFFARX1_RVT PhyAddrPointer_reg_25_ ( .D(n4533), .CLK(CK), .RSTB(n5221), .Q(
        n5081) );
  DFFARX1_RVT rEIP_reg_25_ ( .D(n4595), .CLK(CK), .RSTB(n5221), .Q(rEIP[25])
         );
  DFFARX1_RVT InstAddrPointer_reg_25_ ( .D(n4747), .CLK(CK), .RSTB(n5248), .Q(
        n4917) );
  DFFARX1_RVT PhyAddrPointer_reg_26_ ( .D(n4532), .CLK(CK), .RSTB(n5221), .Q(
        n5082) );
  DFFARX1_RVT rEIP_reg_26_ ( .D(n4594), .CLK(CK), .RSTB(n5221), .Q(rEIP[26])
         );
  DFFARX1_RVT InstAddrPointer_reg_26_ ( .D(n4748), .CLK(CK), .RSTB(n5248), .Q(
        n4979), .QN(n9571) );
  DFFARX1_RVT PhyAddrPointer_reg_27_ ( .D(n4531), .CLK(CK), .RSTB(n5220), .Q(
        n5083) );
  DFFARX1_RVT rEIP_reg_27_ ( .D(n4593), .CLK(CK), .RSTB(n5221), .Q(rEIP[27])
         );
  DFFARX1_RVT InstAddrPointer_reg_27_ ( .D(n4749), .CLK(CK), .RSTB(n5247), .Q(
        n4916) );
  DFFARX1_RVT PhyAddrPointer_reg_28_ ( .D(n4530), .CLK(CK), .RSTB(n5220), .Q(
        n5084) );
  DFFARX1_RVT rEIP_reg_28_ ( .D(n4592), .CLK(CK), .RSTB(n5220), .Q(rEIP[28])
         );
  DFFARX1_RVT InstAddrPointer_reg_28_ ( .D(n4750), .CLK(CK), .RSTB(n5247), .Q(
        n4970), .QN(n9570) );
  DFFARX1_RVT PhyAddrPointer_reg_29_ ( .D(n4529), .CLK(CK), .RSTB(n5220), .Q(
        n5085) );
  DFFARX1_RVT rEIP_reg_29_ ( .D(n4591), .CLK(CK), .RSTB(n5220), .Q(rEIP[29])
         );
  DFFARX1_RVT Address_reg_0_ ( .D(n4588), .CLK(CK), .RSTB(n5216), .Q(
        Address[0]) );
  DFFARX1_RVT Address_reg_1_ ( .D(n4587), .CLK(CK), .RSTB(n5216), .Q(
        Address[1]) );
  DFFARX1_RVT Address_reg_2_ ( .D(n4586), .CLK(CK), .RSTB(n5216), .Q(
        Address[2]) );
  DFFARX1_RVT Address_reg_3_ ( .D(n4585), .CLK(CK), .RSTB(n5216), .Q(
        Address[3]) );
  DFFARX1_RVT Address_reg_4_ ( .D(n4584), .CLK(CK), .RSTB(n5216), .Q(
        Address[4]) );
  DFFARX1_RVT Address_reg_5_ ( .D(n4583), .CLK(CK), .RSTB(n5216), .Q(
        Address[5]) );
  DFFARX1_RVT Address_reg_6_ ( .D(n4582), .CLK(CK), .RSTB(n5216), .Q(
        Address[6]) );
  DFFARX1_RVT Address_reg_7_ ( .D(n4581), .CLK(CK), .RSTB(n5216), .Q(
        Address[7]) );
  DFFARX1_RVT Address_reg_8_ ( .D(n4580), .CLK(CK), .RSTB(n5216), .Q(
        Address[8]) );
  DFFARX1_RVT Address_reg_9_ ( .D(n4579), .CLK(CK), .RSTB(n5216), .Q(
        Address[9]) );
  DFFARX1_RVT Address_reg_10_ ( .D(n4578), .CLK(CK), .RSTB(n5217), .Q(
        Address[10]) );
  DFFARX1_RVT Address_reg_11_ ( .D(n4577), .CLK(CK), .RSTB(n5217), .Q(
        Address[11]) );
  DFFARX1_RVT Address_reg_12_ ( .D(n4576), .CLK(CK), .RSTB(n5217), .Q(
        Address[12]) );
  DFFARX1_RVT Address_reg_13_ ( .D(n4575), .CLK(CK), .RSTB(n5217), .Q(
        Address[13]) );
  DFFARX1_RVT Address_reg_14_ ( .D(n4574), .CLK(CK), .RSTB(n5217), .Q(
        Address[14]) );
  DFFARX1_RVT Address_reg_15_ ( .D(n4573), .CLK(CK), .RSTB(n5217), .Q(
        Address[15]) );
  DFFARX1_RVT Address_reg_16_ ( .D(n4572), .CLK(CK), .RSTB(n5217), .Q(
        Address[16]) );
  DFFARX1_RVT Address_reg_17_ ( .D(n4571), .CLK(CK), .RSTB(n5217), .Q(
        Address[17]) );
  DFFARX1_RVT Address_reg_18_ ( .D(n4570), .CLK(CK), .RSTB(n5217), .Q(
        Address[18]) );
  DFFARX1_RVT Address_reg_19_ ( .D(n4569), .CLK(CK), .RSTB(n5217), .Q(
        Address[19]) );
  DFFARX1_RVT Address_reg_20_ ( .D(n4568), .CLK(CK), .RSTB(n5217), .Q(
        Address[20]) );
  DFFARX1_RVT Address_reg_21_ ( .D(n4567), .CLK(CK), .RSTB(n5217), .Q(
        Address[21]) );
  DFFARX1_RVT Address_reg_22_ ( .D(n4566), .CLK(CK), .RSTB(n5218), .Q(
        Address[22]) );
  DFFARX1_RVT Address_reg_23_ ( .D(n4565), .CLK(CK), .RSTB(n5218), .Q(
        Address[23]) );
  DFFARX1_RVT Address_reg_24_ ( .D(n4564), .CLK(CK), .RSTB(n5218), .Q(
        Address[24]) );
  DFFARX1_RVT Address_reg_25_ ( .D(n4563), .CLK(CK), .RSTB(n5218), .Q(
        Address[25]) );
  DFFARX1_RVT Address_reg_26_ ( .D(n4562), .CLK(CK), .RSTB(n5218), .Q(
        Address[26]) );
  DFFARX1_RVT Address_reg_27_ ( .D(n4561), .CLK(CK), .RSTB(n5218), .Q(
        Address[27]) );
  DFFARX1_RVT Address_reg_28_ ( .D(n4560), .CLK(CK), .RSTB(n5216), .Q(
        Address[28]) );
  DFFARX1_RVT Address_reg_29_ ( .D(n4559), .CLK(CK), .RSTB(n5216), .Q(
        Address[29]) );
  DFFARX1_RVT InstAddrPointer_reg_29_ ( .D(n4751), .CLK(CK), .RSTB(n5247), .Q(
        n4915) );
  DFFARX1_RVT PhyAddrPointer_reg_30_ ( .D(n4528), .CLK(CK), .RSTB(n5219), .Q(
        n5056) );
  DFFARX1_RVT Datao_reg_30_ ( .D(n4496), .CLK(CK), .RSTB(n5220), .Q(Datao[30])
         );
  DFFARX1_RVT DataWidth_reg_0_ ( .D(n4898), .CLK(CK), .RSTB(n5250), .Q(n4914)
         );
  DFFARX1_RVT DataWidth_reg_1_ ( .D(n4897), .CLK(CK), .RSTB(n5250), .Q(n4968), 
        .QN(n9514) );
  DFFARX1_RVT ByteEnable_reg_3_ ( .D(n4495), .CLK(CK), .RSTB(n5218), .Q(n5190)
         );
  DFFARX1_RVT BE_n_reg_3_ ( .D(n4494), .CLK(CK), .RSTB(n5218), .Q(BE_n[3]) );
  DFFARX1_RVT ByteEnable_reg_2_ ( .D(n4493), .CLK(CK), .RSTB(n5219), .Q(n5191)
         );
  DFFARX1_RVT BE_n_reg_2_ ( .D(n4492), .CLK(CK), .RSTB(n5219), .Q(BE_n[2]) );
  DFFARX1_RVT ByteEnable_reg_1_ ( .D(n4491), .CLK(CK), .RSTB(n5218), .Q(n5192)
         );
  DFFARX1_RVT BE_n_reg_1_ ( .D(n4490), .CLK(CK), .RSTB(n5218), .Q(BE_n[1]) );
  DFFARX1_RVT ByteEnable_reg_0_ ( .D(n4489), .CLK(CK), .RSTB(n5218), .Q(n5193)
         );
  DFFARX1_RVT BE_n_reg_0_ ( .D(n4488), .CLK(CK), .RSTB(n5218), .Q(BE_n[0]) );
  DFFARX2_RVT InstQueueRd_Addr_reg_3_ ( .D(n4760), .CLK(CK), .RSTB(n5246), .Q(
        n4906), .QN(n936) );
  INVX2_RVT U4487 ( .A(n9478), .Y(n9278) );
  NAND3X0_RVT U4488 ( .A1(n9280), .A2(n9281), .A3(n9279), .Y(n9276) );
  INVX2_RVT U4489 ( .A(n6487), .Y(n6516) );
  NAND3X0_RVT U4490 ( .A1(n7871), .A2(n5265), .A3(n8881), .Y(n6445) );
  NAND4X0_RVT U4491 ( .A1(n6446), .A2(n6531), .A3(n6433), .A4(n6755), .Y(n7865) );
  AND2X2_RVT U4492 ( .A1(n7192), .A2(n7052), .Y(n7057) );
  NAND2X0_RVT U4493 ( .A1(n7004), .A2(n5209), .Y(n4963) );
  INVX0_RVT U4494 ( .A(n4963), .Y(n5196) );
  INVX0_RVT U4495 ( .A(n4963), .Y(n5197) );
  INVX0_RVT U4496 ( .A(n4963), .Y(n5198) );
  INVX0_RVT U4497 ( .A(n4963), .Y(n5199) );
  INVX0_RVT U4498 ( .A(n6768), .Y(n5200) );
  INVX0_RVT U4499 ( .A(n6768), .Y(n5201) );
  INVX0_RVT U4500 ( .A(n6768), .Y(n5202) );
  INVX0_RVT U4501 ( .A(n6768), .Y(n5203) );
  INVX0_RVT U4502 ( .A(n7006), .Y(n5204) );
  INVX0_RVT U4503 ( .A(n7006), .Y(n5205) );
  INVX0_RVT U4504 ( .A(n7006), .Y(n5206) );
  INVX0_RVT U4505 ( .A(n7006), .Y(n5207) );
  INVX0_RVT U4506 ( .A(n5200), .Y(n5208) );
  INVX0_RVT U4507 ( .A(n5201), .Y(n5209) );
  INVX0_RVT U4508 ( .A(n5202), .Y(n5210) );
  INVX0_RVT U4509 ( .A(n5203), .Y(n5211) );
  INVX0_RVT U4510 ( .A(n6432), .Y(n5212) );
  INVX0_RVT U4511 ( .A(n6432), .Y(n5213) );
  INVX0_RVT U4512 ( .A(n6432), .Y(n5214) );
  INVX0_RVT U4513 ( .A(n6432), .Y(n5215) );
  INVX2_RVT U4514 ( .A(n8507), .Y(n8881) );
  AND3X2_RVT U4515 ( .A1(n6321), .A2(n6330), .A3(n7844), .Y(n7192) );
  AND2X2_RVT U4516 ( .A1(n938), .A2(n939), .Y(n7842) );
  NAND3X2_RVT U4517 ( .A1(n6380), .A2(n6381), .A3(n6382), .Y(n5330) );
  AND2X2_RVT U4518 ( .A1(n939), .A2(n4927), .Y(n7852) );
  AND2X2_RVT U4519 ( .A1(n5265), .A2(n8673), .Y(n8565) );
  AND2X2_RVT U4520 ( .A1(n5265), .A2(n8558), .Y(n8110) );
  AND2X1_RVT U4521 ( .A1(n5265), .A2(n5323), .Y(n6725) );
  INVX2_RVT U4522 ( .A(n6407), .Y(n5265) );
  XOR2X2_RVT U4523 ( .A1(n7259), .A2(n6377), .Y(n5431) );
  AND2X2_RVT U4524 ( .A1(n4927), .A2(n4908), .Y(n7848) );
  INVX2_RVT U4525 ( .A(n5363), .Y(n5359) );
  INVX2_RVT U4526 ( .A(n6433), .Y(n8114) );
  NAND2X2_RVT U4527 ( .A1(n8560), .A2(n6760), .Y(n6433) );
  NAND2X2_RVT U4528 ( .A1(n7007), .A2(n7197), .Y(n7430) );
  INVX2_RVT U4529 ( .A(n7045), .Y(n6863) );
  NAND2X2_RVT U4530 ( .A1(n8950), .A2(n5390), .Y(n8108) );
  AND2X2_RVT U4531 ( .A1(n7207), .A2(n7866), .Y(n7212) );
  INVX4_RVT U4532 ( .A(n8192), .Y(n8112) );
  INVX4_RVT U4533 ( .A(n5351), .Y(n5371) );
  NAND2X4_RVT U4534 ( .A1(n7908), .A2(n6422), .Y(n7217) );
  AND2X4_RVT U4535 ( .A1(n936), .A2(n937), .Y(n7694) );
  AND2X2_RVT U4536 ( .A1(n938), .A2(n4908), .Y(n7853) );
  INVX2_RVT U4537 ( .A(n5390), .Y(n5476) );
  INVX2_RVT U4538 ( .A(n5323), .Y(n6545) );
  INVX2_RVT U4539 ( .A(n5279), .Y(n8035) );
  NAND2X2_RVT U4540 ( .A1(n7862), .A2(n7863), .Y(n7214) );
  AND3X2_RVT U4541 ( .A1(n6422), .A2(n7869), .A3(n7207), .Y(n7210) );
  AND2X2_RVT U4542 ( .A1(n5272), .A2(n7045), .Y(n6864) );
  INVX2_RVT U4543 ( .A(n8673), .Y(n8568) );
  INVX2_RVT U4544 ( .A(n5301), .Y(n8036) );
  AND2X2_RVT U4545 ( .A1(n6725), .A2(n6726), .Y(n5319) );
  AND2X2_RVT U4546 ( .A1(n6725), .A2(n6730), .Y(n5321) );
  NAND2X2_RVT U4547 ( .A1(n6445), .A2(n9160), .Y(n8109) );
  INVX2_RVT U4548 ( .A(n8558), .Y(n8113) );
  INVX2_RVT U4549 ( .A(n6446), .Y(n7215) );
  INVX2_RVT U4550 ( .A(n7865), .Y(n7218) );
  INVX2_RVT U4551 ( .A(n7052), .Y(n7051) );
  NAND2X4_RVT U4552 ( .A1(n7197), .A2(n7198), .Y(n7052) );
  INVX4_RVT U4553 ( .A(n6751), .Y(n5276) );
  INVX2_RVT U4554 ( .A(n6422), .Y(n7864) );
  NAND3X4_RVT U4555 ( .A1(n8927), .A2(n8928), .A3(n8929), .Y(n6422) );
  NAND2X4_RVT U4556 ( .A1(n5351), .A2(n5368), .Y(n5479) );
  AND2X4_RVT U4557 ( .A1(n937), .A2(n4906), .Y(n7766) );
  NAND2X4_RVT U4558 ( .A1(n8515), .A2(n6739), .Y(n8192) );
  AND2X4_RVT U4559 ( .A1(n936), .A2(n4926), .Y(n7678) );
  NBUFFX4_RVT U4560 ( .A(n9581), .Y(n5254) );
  NBUFFX4_RVT U4561 ( .A(n9581), .Y(n5252) );
  NBUFFX4_RVT U4562 ( .A(n9581), .Y(n5253) );
  NBUFFX4_RVT U4563 ( .A(n9581), .Y(n5255) );
  NBUFFX4_RVT U4564 ( .A(n9581), .Y(n5251) );
  NBUFFX4_RVT U4565 ( .A(n5255), .Y(n5216) );
  NBUFFX4_RVT U4566 ( .A(n5255), .Y(n5217) );
  NBUFFX4_RVT U4567 ( .A(n5255), .Y(n5218) );
  NBUFFX4_RVT U4568 ( .A(n5255), .Y(n5219) );
  NBUFFX4_RVT U4569 ( .A(n5255), .Y(n5220) );
  NBUFFX4_RVT U4570 ( .A(n5255), .Y(n5221) );
  NBUFFX4_RVT U4571 ( .A(n5255), .Y(n5222) );
  NBUFFX4_RVT U4572 ( .A(n5254), .Y(n5223) );
  NBUFFX4_RVT U4573 ( .A(n5254), .Y(n5224) );
  NBUFFX4_RVT U4574 ( .A(n5254), .Y(n5225) );
  NBUFFX4_RVT U4575 ( .A(n5254), .Y(n5226) );
  NBUFFX4_RVT U4576 ( .A(n5254), .Y(n5227) );
  NBUFFX4_RVT U4577 ( .A(n5254), .Y(n5228) );
  NBUFFX4_RVT U4578 ( .A(n5254), .Y(n5229) );
  NBUFFX4_RVT U4579 ( .A(n5253), .Y(n5230) );
  NBUFFX4_RVT U4580 ( .A(n5253), .Y(n5231) );
  NBUFFX4_RVT U4581 ( .A(n5253), .Y(n5232) );
  NBUFFX4_RVT U4582 ( .A(n5253), .Y(n5233) );
  NBUFFX4_RVT U4583 ( .A(n5253), .Y(n5234) );
  NBUFFX4_RVT U4584 ( .A(n5253), .Y(n5235) );
  NBUFFX4_RVT U4585 ( .A(n5253), .Y(n5236) );
  NBUFFX4_RVT U4586 ( .A(n5252), .Y(n5237) );
  NBUFFX4_RVT U4587 ( .A(n5252), .Y(n5238) );
  NBUFFX4_RVT U4588 ( .A(n5252), .Y(n5239) );
  NBUFFX4_RVT U4589 ( .A(n5252), .Y(n5240) );
  NBUFFX4_RVT U4590 ( .A(n5252), .Y(n5241) );
  NBUFFX4_RVT U4591 ( .A(n5252), .Y(n5242) );
  NBUFFX4_RVT U4592 ( .A(n5252), .Y(n5243) );
  NBUFFX4_RVT U4593 ( .A(n5251), .Y(n5244) );
  NBUFFX4_RVT U4594 ( .A(n5251), .Y(n5245) );
  NBUFFX4_RVT U4595 ( .A(n5251), .Y(n5246) );
  NBUFFX4_RVT U4596 ( .A(n5251), .Y(n5247) );
  NBUFFX4_RVT U4597 ( .A(n5251), .Y(n5248) );
  NBUFFX4_RVT U4598 ( .A(n5251), .Y(n5249) );
  NBUFFX4_RVT U4599 ( .A(n5251), .Y(n5250) );
  INVX0_RVT U4600 ( .A(reset), .Y(n9581) );
  NAND2X0_RVT U4601 ( .A1(n5256), .A2(n5257), .Y(n4904) );
  OR2X1_RVT U4602 ( .A1(n5258), .A2(n979), .Y(n5257) );
  NAND2X0_RVT U4603 ( .A1(n5259), .A2(n5258), .Y(n5256) );
  NAND2X0_RVT U4604 ( .A1(n5260), .A2(n5261), .Y(n5258) );
  NAND3X0_RVT U4605 ( .A1(n5262), .A2(n5263), .A3(n5264), .Y(n5259) );
  NAND2X0_RVT U4606 ( .A1(n5265), .A2(n5266), .Y(n5262) );
  NAND3X0_RVT U4607 ( .A1(n5267), .A2(n5268), .A3(n5269), .Y(n5266) );
  OR2X1_RVT U4608 ( .A1(n5270), .A2(n5271), .Y(n5269) );
  NAND2X0_RVT U4609 ( .A1(n5272), .A2(n5273), .Y(n5267) );
  NAND2X0_RVT U4610 ( .A1(n4967), .A2(n5271), .Y(n5273) );
  AND2X1_RVT U4611 ( .A1(n5274), .A2(n5275), .Y(n4903) );
  NAND3X0_RVT U4612 ( .A1(n5276), .A2(n5277), .A3(NA_n), .Y(n5275) );
  NAND2X0_RVT U4613 ( .A1(n5278), .A2(n4929), .Y(n5277) );
  NAND4X0_RVT U4614 ( .A1(n5279), .A2(n5280), .A3(n5281), .A4(n5282), .Y(n5274) );
  AND2X1_RVT U4615 ( .A1(n5283), .A2(n5284), .Y(n5282) );
  NAND4X0_RVT U4616 ( .A1(n979), .A2(HOLD), .A3(n731), .A4(n4929), .Y(n5284)
         );
  NAND2X0_RVT U4617 ( .A1(READY_n), .A2(n5285), .Y(n5283) );
  NAND2X0_RVT U4618 ( .A1(n5286), .A2(n5287), .Y(n5285) );
  NAND2X0_RVT U4619 ( .A1(n5288), .A2(n5289), .Y(n5287) );
  NAND2X0_RVT U4620 ( .A1(n979), .A2(n5290), .Y(n5289) );
  INVX0_RVT U4621 ( .A(n5291), .Y(n5288) );
  NAND2X0_RVT U4622 ( .A1(n4913), .A2(n4962), .Y(n5286) );
  NAND4X0_RVT U4623 ( .A1(n5292), .A2(n5293), .A3(n5294), .A4(n5291), .Y(n4902) );
  NAND3X0_RVT U4624 ( .A1(n5295), .A2(n4929), .A3(n5296), .Y(n5291) );
  NAND2X0_RVT U4625 ( .A1(n5290), .A2(n5268), .Y(n5295) );
  NAND2X0_RVT U4626 ( .A1(n5297), .A2(n4929), .Y(n5292) );
  NAND4X0_RVT U4627 ( .A1(n5298), .A2(n5299), .A3(n5293), .A4(n5280), .Y(n4901) );
  NAND2X0_RVT U4628 ( .A1(n5271), .A2(n5300), .Y(n5293) );
  NAND4X0_RVT U4629 ( .A1(n5301), .A2(n5290), .A3(n5302), .A4(n4989), .Y(n5300) );
  INVX0_RVT U4630 ( .A(NA_n), .Y(n5302) );
  INVX0_RVT U4631 ( .A(HOLD), .Y(n5290) );
  NAND2X0_RVT U4632 ( .A1(READY_n), .A2(n4962), .Y(n5299) );
  NAND2X0_RVT U4633 ( .A1(n5303), .A2(n4929), .Y(n5298) );
  NAND2X0_RVT U4634 ( .A1(n5304), .A2(n5297), .Y(n5303) );
  NAND2X0_RVT U4635 ( .A1(n5281), .A2(n4989), .Y(n5297) );
  NAND2X0_RVT U4636 ( .A1(HOLD), .A2(n4913), .Y(n5281) );
  NAND2X0_RVT U4637 ( .A1(HOLD), .A2(n5296), .Y(n5304) );
  NAND3X0_RVT U4638 ( .A1(n5305), .A2(n5294), .A3(n5306), .Y(n4900) );
  NAND2X0_RVT U4639 ( .A1(n5276), .A2(ADS_n), .Y(n5305) );
  NAND2X0_RVT U4640 ( .A1(n5307), .A2(n5308), .Y(n4899) );
  NAND2X0_RVT U4641 ( .A1(n5306), .A2(n4967), .Y(n5308) );
  NAND2X0_RVT U4642 ( .A1(n5309), .A2(n5310), .Y(n4898) );
  OR2X1_RVT U4643 ( .A1(n5306), .A2(BS16_n), .Y(n5310) );
  NAND3X0_RVT U4644 ( .A1(n5294), .A2(n4914), .A3(n5306), .Y(n5309) );
  NAND2X0_RVT U4645 ( .A1(n5307), .A2(n5311), .Y(n4897) );
  NAND2X0_RVT U4646 ( .A1(n5306), .A2(n4968), .Y(n5311) );
  INVX0_RVT U4647 ( .A(n5312), .Y(n5306) );
  AND2X1_RVT U4648 ( .A1(n5294), .A2(n5313), .Y(n5307) );
  NAND2X0_RVT U4649 ( .A1(BS16_n), .A2(n5312), .Y(n5313) );
  NAND2X0_RVT U4650 ( .A1(n5280), .A2(n5314), .Y(n5312) );
  NAND2X0_RVT U4651 ( .A1(n5296), .A2(n4929), .Y(n5314) );
  NAND4X0_RVT U4652 ( .A1(n5315), .A2(n5316), .A3(n5317), .A4(n5318), .Y(n4896) );
  NAND2X0_RVT U4653 ( .A1(n5319), .A2(n5320), .Y(n5318) );
  NAND2X0_RVT U4654 ( .A1(n5321), .A2(n5322), .Y(n5317) );
  OR2X1_RVT U4655 ( .A1(n5323), .A2(n9567), .Y(n5316) );
  NAND3X0_RVT U4656 ( .A1(n5325), .A2(n5326), .A3(n5327), .Y(n4894) );
  NAND2X0_RVT U4657 ( .A1(n5328), .A2(n5329), .Y(n5327) );
  OR2X1_RVT U4658 ( .A1(n5330), .A2(n801), .Y(n5326) );
  NAND2X0_RVT U4659 ( .A1(n5331), .A2(n5330), .Y(n5325) );
  NAND3X0_RVT U4660 ( .A1(n5332), .A2(n5333), .A3(n5334), .Y(n5331) );
  NAND2X0_RVT U4661 ( .A1(n5335), .A2(n5336), .Y(n5333) );
  NAND2X0_RVT U4662 ( .A1(n5337), .A2(n5338), .Y(n5332) );
  NAND3X0_RVT U4663 ( .A1(n5339), .A2(n5340), .A3(n5341), .Y(n4893) );
  NAND2X0_RVT U4664 ( .A1(n5342), .A2(n4925), .Y(n5341) );
  NAND2X0_RVT U4665 ( .A1(n5343), .A2(n5344), .Y(n4892) );
  NAND2X0_RVT U4666 ( .A1(n5345), .A2(n5346), .Y(n5344) );
  OR2X1_RVT U4667 ( .A1(n5347), .A2(n974), .Y(n5346) );
  NAND2X0_RVT U4668 ( .A1(n5348), .A2(n4909), .Y(n5343) );
  NAND2X0_RVT U4669 ( .A1(n5349), .A2(n5350), .Y(n5348) );
  OR2X1_RVT U4670 ( .A1(n5345), .A2(n5351), .Y(n5350) );
  XOR2X1_RVT U4671 ( .A1(n5352), .A2(n5353), .Y(n5345) );
  NAND3X0_RVT U4672 ( .A1(n5354), .A2(n5355), .A3(n5356), .Y(n4891) );
  NAND3X0_RVT U4673 ( .A1(n5357), .A2(n5349), .A3(n5358), .Y(n5356) );
  NAND2X0_RVT U4674 ( .A1(n5359), .A2(n975), .Y(n5355) );
  NAND2X0_RVT U4675 ( .A1(n5360), .A2(n4928), .Y(n5354) );
  NAND3X0_RVT U4676 ( .A1(n5349), .A2(n5351), .A3(n5361), .Y(n5360) );
  NAND2X0_RVT U4677 ( .A1(n5362), .A2(n5363), .Y(n5361) );
  NAND3X0_RVT U4678 ( .A1(n5364), .A2(n5365), .A3(n5366), .Y(n4890) );
  NAND2X0_RVT U4679 ( .A1(n5367), .A2(n5347), .Y(n5366) );
  NAND2X0_RVT U4680 ( .A1(n5340), .A2(n5368), .Y(n5347) );
  INVX0_RVT U4681 ( .A(n5369), .Y(n5367) );
  NAND2X0_RVT U4682 ( .A1(n5370), .A2(n4907), .Y(n5365) );
  NAND3X0_RVT U4683 ( .A1(n5371), .A2(n5372), .A3(n973), .Y(n5364) );
  NAND2X0_RVT U4684 ( .A1(n5373), .A2(n5374), .Y(n4889) );
  NAND2X0_RVT U4685 ( .A1(n5375), .A2(n4930), .Y(n5374) );
  NAND3X0_RVT U4686 ( .A1(n5376), .A2(n5377), .A3(n5378), .Y(n5375) );
  INVX0_RVT U4687 ( .A(n5370), .Y(n5378) );
  NAND2X0_RVT U4688 ( .A1(n5349), .A2(n5379), .Y(n5370) );
  OR2X1_RVT U4689 ( .A1(n5372), .A2(n5351), .Y(n5379) );
  NAND4X0_RVT U4690 ( .A1(n5380), .A2(n5381), .A3(n5363), .A4(n5382), .Y(n5349) );
  NAND2X0_RVT U4691 ( .A1(n5357), .A2(n5383), .Y(n5381) );
  NAND2X0_RVT U4692 ( .A1(n5384), .A2(n5362), .Y(n5377) );
  NAND2X0_RVT U4693 ( .A1(n5371), .A2(n973), .Y(n5376) );
  NAND2X0_RVT U4694 ( .A1(n965), .A2(n5385), .Y(n5373) );
  NAND2X0_RVT U4695 ( .A1(n5384), .A2(n5386), .Y(n5385) );
  NAND3X0_RVT U4696 ( .A1(n5372), .A2(n4907), .A3(n5371), .Y(n5386) );
  NAND2X0_RVT U4697 ( .A1(n974), .A2(n5369), .Y(n5372) );
  NAND2X0_RVT U4698 ( .A1(n5384), .A2(n5387), .Y(n5369) );
  NAND2X0_RVT U4699 ( .A1(n5388), .A2(n5389), .Y(n5387) );
  OR2X1_RVT U4700 ( .A1(n5389), .A2(n5388), .Y(n5384) );
  NAND2X0_RVT U4701 ( .A1(n4907), .A2(n5362), .Y(n5388) );
  NAND2X0_RVT U4702 ( .A1(n5352), .A2(n5353), .Y(n5389) );
  NAND2X0_RVT U4703 ( .A1(n5390), .A2(n5391), .Y(n5353) );
  NAND2X0_RVT U4704 ( .A1(n5362), .A2(n4909), .Y(n5391) );
  NAND2X0_RVT U4705 ( .A1(n5368), .A2(n5363), .Y(n5362) );
  NAND2X0_RVT U4706 ( .A1(n5380), .A2(n5392), .Y(n5352) );
  NAND2X0_RVT U4707 ( .A1(n5359), .A2(n4928), .Y(n5392) );
  NAND3X0_RVT U4708 ( .A1(n5393), .A2(n5394), .A3(n5395), .Y(n4888) );
  NAND2X0_RVT U4709 ( .A1(n5396), .A2(n5397), .Y(n5395) );
  NAND2X0_RVT U4710 ( .A1(n5398), .A2(n5118), .Y(n5394) );
  NAND2X0_RVT U4711 ( .A1(n5399), .A2(n5400), .Y(n5393) );
  NAND3X0_RVT U4712 ( .A1(n5401), .A2(n5402), .A3(n5403), .Y(n5399) );
  NAND2X0_RVT U4713 ( .A1(n5404), .A2(n5405), .Y(n5402) );
  NAND2X0_RVT U4714 ( .A1(n5406), .A2(n5407), .Y(n5401) );
  NAND3X0_RVT U4715 ( .A1(n5408), .A2(n5409), .A3(n5410), .Y(n4887) );
  NAND2X0_RVT U4716 ( .A1(n5396), .A2(n5411), .Y(n5410) );
  NAND2X0_RVT U4717 ( .A1(n5398), .A2(n5128), .Y(n5409) );
  NAND2X0_RVT U4718 ( .A1(n5412), .A2(n5400), .Y(n5408) );
  NAND3X0_RVT U4719 ( .A1(n5413), .A2(n5414), .A3(n5415), .Y(n5412) );
  NAND2X0_RVT U4720 ( .A1(n5416), .A2(n5405), .Y(n5414) );
  NAND2X0_RVT U4721 ( .A1(n5406), .A2(n5417), .Y(n5413) );
  NAND3X0_RVT U4722 ( .A1(n5418), .A2(n5419), .A3(n5420), .Y(n4886) );
  NAND2X0_RVT U4723 ( .A1(n5421), .A2(n5396), .Y(n5420) );
  NAND2X0_RVT U4724 ( .A1(n5398), .A2(n5131), .Y(n5419) );
  NAND2X0_RVT U4725 ( .A1(n5422), .A2(n5400), .Y(n5418) );
  NAND3X0_RVT U4726 ( .A1(n5423), .A2(n5424), .A3(n5425), .Y(n5422) );
  NAND2X0_RVT U4727 ( .A1(n5426), .A2(n5405), .Y(n5424) );
  NAND2X0_RVT U4728 ( .A1(n5406), .A2(n5427), .Y(n5423) );
  NAND3X0_RVT U4729 ( .A1(n5428), .A2(n5429), .A3(n5430), .Y(n4885) );
  NAND2X0_RVT U4730 ( .A1(n5431), .A2(n5396), .Y(n5430) );
  NAND2X0_RVT U4731 ( .A1(n5398), .A2(n5119), .Y(n5429) );
  NAND2X0_RVT U4732 ( .A1(n5432), .A2(n5400), .Y(n5428) );
  NAND3X0_RVT U4733 ( .A1(n5433), .A2(n5434), .A3(n5435), .Y(n5432) );
  NAND2X0_RVT U4734 ( .A1(n5436), .A2(n5405), .Y(n5434) );
  NAND2X0_RVT U4735 ( .A1(n5406), .A2(n5437), .Y(n5433) );
  NAND3X0_RVT U4736 ( .A1(n5438), .A2(n5439), .A3(n5440), .Y(n4884) );
  NAND2X0_RVT U4737 ( .A1(n5441), .A2(n5396), .Y(n5440) );
  NAND2X0_RVT U4738 ( .A1(n5398), .A2(n5120), .Y(n5439) );
  NAND2X0_RVT U4739 ( .A1(n5442), .A2(n5400), .Y(n5438) );
  NAND3X0_RVT U4740 ( .A1(n5443), .A2(n5444), .A3(n5445), .Y(n5442) );
  NAND2X0_RVT U4741 ( .A1(n5446), .A2(n5405), .Y(n5444) );
  NAND2X0_RVT U4742 ( .A1(n5447), .A2(n5406), .Y(n5443) );
  NAND3X0_RVT U4743 ( .A1(n5448), .A2(n5449), .A3(n5450), .Y(n4883) );
  NAND2X0_RVT U4744 ( .A1(n5451), .A2(n5396), .Y(n5450) );
  NAND2X0_RVT U4745 ( .A1(n5398), .A2(n5121), .Y(n5449) );
  NAND2X0_RVT U4746 ( .A1(n5452), .A2(n5400), .Y(n5448) );
  NAND3X0_RVT U4747 ( .A1(n5453), .A2(n5454), .A3(n5455), .Y(n5452) );
  NAND2X0_RVT U4748 ( .A1(n5456), .A2(n5405), .Y(n5454) );
  NAND2X0_RVT U4749 ( .A1(n5406), .A2(n5457), .Y(n5453) );
  NAND3X0_RVT U4750 ( .A1(n5458), .A2(n5459), .A3(n5460), .Y(n4882) );
  NAND2X0_RVT U4751 ( .A1(n5396), .A2(n5461), .Y(n5460) );
  NAND2X0_RVT U4752 ( .A1(n5398), .A2(n5122), .Y(n5459) );
  NAND2X0_RVT U4753 ( .A1(n5462), .A2(n5400), .Y(n5458) );
  NAND3X0_RVT U4754 ( .A1(n5463), .A2(n5464), .A3(n5465), .Y(n5462) );
  NAND2X0_RVT U4755 ( .A1(n5466), .A2(n5405), .Y(n5464) );
  NAND2X0_RVT U4756 ( .A1(n5406), .A2(n5467), .Y(n5463) );
  NAND3X0_RVT U4757 ( .A1(n5468), .A2(n5469), .A3(n5470), .Y(n4881) );
  NAND2X0_RVT U4758 ( .A1(n5396), .A2(n5329), .Y(n5470) );
  AND2X1_RVT U4759 ( .A1(n5471), .A2(n5400), .Y(n5396) );
  NAND2X0_RVT U4760 ( .A1(n5398), .A2(n5049), .Y(n5469) );
  INVX0_RVT U4761 ( .A(n5400), .Y(n5398) );
  NAND2X0_RVT U4762 ( .A1(n5472), .A2(n5400), .Y(n5468) );
  NAND3X0_RVT U4763 ( .A1(n5473), .A2(n5474), .A3(n5475), .Y(n5400) );
  NAND2X0_RVT U4764 ( .A1(n5476), .A2(n5477), .Y(n5475) );
  NAND2X0_RVT U4765 ( .A1(n5478), .A2(n5479), .Y(n5474) );
  NAND2X0_RVT U4766 ( .A1(n5480), .A2(n5359), .Y(n5473) );
  NAND3X0_RVT U4767 ( .A1(n5481), .A2(n5482), .A3(n5334), .Y(n5472) );
  NAND2X0_RVT U4768 ( .A1(n5405), .A2(n5335), .Y(n5482) );
  INVX0_RVT U4769 ( .A(n5477), .Y(n5405) );
  NAND2X0_RVT U4770 ( .A1(n5338), .A2(n5406), .Y(n5481) );
  NAND3X0_RVT U4771 ( .A1(n5483), .A2(n5484), .A3(n5485), .Y(n4880) );
  NAND2X0_RVT U4772 ( .A1(n5486), .A2(n5397), .Y(n5485) );
  NAND2X0_RVT U4773 ( .A1(n5487), .A2(n5123), .Y(n5484) );
  NAND2X0_RVT U4774 ( .A1(n5488), .A2(n5489), .Y(n5483) );
  NAND3X0_RVT U4775 ( .A1(n5490), .A2(n5491), .A3(n5403), .Y(n5488) );
  NAND2X0_RVT U4776 ( .A1(n5492), .A2(n5404), .Y(n5491) );
  NAND2X0_RVT U4777 ( .A1(n5471), .A2(n5407), .Y(n5490) );
  NAND3X0_RVT U4778 ( .A1(n5493), .A2(n5494), .A3(n5495), .Y(n4879) );
  NAND2X0_RVT U4779 ( .A1(n5486), .A2(n5411), .Y(n5495) );
  NAND2X0_RVT U4780 ( .A1(n5487), .A2(n5129), .Y(n5494) );
  NAND2X0_RVT U4781 ( .A1(n5496), .A2(n5489), .Y(n5493) );
  NAND3X0_RVT U4782 ( .A1(n5497), .A2(n5498), .A3(n5415), .Y(n5496) );
  NAND2X0_RVT U4783 ( .A1(n5492), .A2(n5416), .Y(n5498) );
  NAND2X0_RVT U4784 ( .A1(n5471), .A2(n5417), .Y(n5497) );
  NAND3X0_RVT U4785 ( .A1(n5499), .A2(n5500), .A3(n5501), .Y(n4878) );
  NAND2X0_RVT U4786 ( .A1(n5486), .A2(n5421), .Y(n5501) );
  NAND2X0_RVT U4787 ( .A1(n5487), .A2(n5130), .Y(n5500) );
  NAND2X0_RVT U4788 ( .A1(n5502), .A2(n5489), .Y(n5499) );
  NAND3X0_RVT U4789 ( .A1(n5503), .A2(n5504), .A3(n5425), .Y(n5502) );
  NAND2X0_RVT U4790 ( .A1(n5492), .A2(n5426), .Y(n5504) );
  NAND2X0_RVT U4791 ( .A1(n5471), .A2(n5427), .Y(n5503) );
  NAND3X0_RVT U4792 ( .A1(n5505), .A2(n5506), .A3(n5507), .Y(n4877) );
  NAND2X0_RVT U4793 ( .A1(n5486), .A2(n5431), .Y(n5507) );
  NAND2X0_RVT U4794 ( .A1(n5487), .A2(n5124), .Y(n5506) );
  NAND2X0_RVT U4795 ( .A1(n5508), .A2(n5489), .Y(n5505) );
  NAND3X0_RVT U4796 ( .A1(n5509), .A2(n5510), .A3(n5435), .Y(n5508) );
  NAND2X0_RVT U4797 ( .A1(n5492), .A2(n5436), .Y(n5510) );
  NAND2X0_RVT U4798 ( .A1(n5471), .A2(n5437), .Y(n5509) );
  NAND3X0_RVT U4799 ( .A1(n5511), .A2(n5512), .A3(n5513), .Y(n4876) );
  NAND2X0_RVT U4800 ( .A1(n5486), .A2(n5441), .Y(n5513) );
  NAND2X0_RVT U4801 ( .A1(n5487), .A2(n5125), .Y(n5512) );
  NAND2X0_RVT U4802 ( .A1(n5514), .A2(n5489), .Y(n5511) );
  NAND3X0_RVT U4803 ( .A1(n5515), .A2(n5516), .A3(n5445), .Y(n5514) );
  NAND2X0_RVT U4804 ( .A1(n5492), .A2(n5446), .Y(n5516) );
  NAND2X0_RVT U4805 ( .A1(n5447), .A2(n5471), .Y(n5515) );
  NAND3X0_RVT U4806 ( .A1(n5517), .A2(n5518), .A3(n5519), .Y(n4875) );
  NAND2X0_RVT U4807 ( .A1(n5486), .A2(n5451), .Y(n5519) );
  NAND2X0_RVT U4808 ( .A1(n5487), .A2(n5126), .Y(n5518) );
  NAND2X0_RVT U4809 ( .A1(n5520), .A2(n5489), .Y(n5517) );
  NAND3X0_RVT U4810 ( .A1(n5521), .A2(n5522), .A3(n5455), .Y(n5520) );
  NAND2X0_RVT U4811 ( .A1(n5492), .A2(n5456), .Y(n5522) );
  NAND2X0_RVT U4812 ( .A1(n5471), .A2(n5457), .Y(n5521) );
  NAND3X0_RVT U4813 ( .A1(n5523), .A2(n5524), .A3(n5525), .Y(n4874) );
  NAND2X0_RVT U4814 ( .A1(n5486), .A2(n5461), .Y(n5525) );
  NAND2X0_RVT U4815 ( .A1(n5487), .A2(n5127), .Y(n5524) );
  NAND2X0_RVT U4816 ( .A1(n5526), .A2(n5489), .Y(n5523) );
  NAND3X0_RVT U4817 ( .A1(n5527), .A2(n5528), .A3(n5465), .Y(n5526) );
  NAND2X0_RVT U4818 ( .A1(n5492), .A2(n5466), .Y(n5528) );
  NAND2X0_RVT U4819 ( .A1(n5471), .A2(n5467), .Y(n5527) );
  NAND3X0_RVT U4820 ( .A1(n5529), .A2(n5530), .A3(n5531), .Y(n4873) );
  NAND2X0_RVT U4821 ( .A1(n5486), .A2(n5329), .Y(n5531) );
  AND2X1_RVT U4822 ( .A1(n5532), .A2(n5489), .Y(n5486) );
  NAND2X0_RVT U4823 ( .A1(n5487), .A2(n5167), .Y(n5530) );
  INVX0_RVT U4824 ( .A(n5489), .Y(n5487) );
  NAND2X0_RVT U4825 ( .A1(n5533), .A2(n5489), .Y(n5529) );
  NAND3X0_RVT U4826 ( .A1(n5534), .A2(n5535), .A3(n5536), .Y(n5489) );
  NAND2X0_RVT U4827 ( .A1(n5476), .A2(n5537), .Y(n5536) );
  NAND2X0_RVT U4828 ( .A1(n5538), .A2(n5479), .Y(n5535) );
  NAND2X0_RVT U4829 ( .A1(n5539), .A2(n5359), .Y(n5534) );
  NAND3X0_RVT U4830 ( .A1(n5540), .A2(n5541), .A3(n5334), .Y(n5533) );
  NAND2X0_RVT U4831 ( .A1(n5492), .A2(n5335), .Y(n5541) );
  INVX0_RVT U4832 ( .A(n5537), .Y(n5492) );
  NAND2X0_RVT U4833 ( .A1(n5471), .A2(n5338), .Y(n5540) );
  NAND3X0_RVT U4834 ( .A1(n5542), .A2(n5543), .A3(n5544), .Y(n4872) );
  NAND2X0_RVT U4835 ( .A1(n5545), .A2(n5397), .Y(n5544) );
  NAND2X0_RVT U4836 ( .A1(n5546), .A2(n5132), .Y(n5543) );
  NAND2X0_RVT U4837 ( .A1(n5547), .A2(n5548), .Y(n5542) );
  NAND3X0_RVT U4838 ( .A1(n5549), .A2(n5550), .A3(n5403), .Y(n5547) );
  NAND2X0_RVT U4839 ( .A1(n5551), .A2(n5404), .Y(n5550) );
  NAND2X0_RVT U4840 ( .A1(n5532), .A2(n5407), .Y(n5549) );
  NAND3X0_RVT U4841 ( .A1(n5552), .A2(n5553), .A3(n5554), .Y(n4871) );
  NAND2X0_RVT U4842 ( .A1(n5545), .A2(n5411), .Y(n5554) );
  NAND2X0_RVT U4843 ( .A1(n5546), .A2(n5137), .Y(n5553) );
  NAND2X0_RVT U4844 ( .A1(n5555), .A2(n5548), .Y(n5552) );
  NAND3X0_RVT U4845 ( .A1(n5556), .A2(n5557), .A3(n5415), .Y(n5555) );
  NAND2X0_RVT U4846 ( .A1(n5551), .A2(n5416), .Y(n5557) );
  NAND2X0_RVT U4847 ( .A1(n5532), .A2(n5417), .Y(n5556) );
  NAND3X0_RVT U4848 ( .A1(n5558), .A2(n5559), .A3(n5560), .Y(n4870) );
  NAND2X0_RVT U4849 ( .A1(n5545), .A2(n5421), .Y(n5560) );
  NAND2X0_RVT U4850 ( .A1(n5546), .A2(n5142), .Y(n5559) );
  NAND2X0_RVT U4851 ( .A1(n5561), .A2(n5548), .Y(n5558) );
  NAND3X0_RVT U4852 ( .A1(n5562), .A2(n5563), .A3(n5425), .Y(n5561) );
  NAND2X0_RVT U4853 ( .A1(n5551), .A2(n5426), .Y(n5563) );
  NAND2X0_RVT U4854 ( .A1(n5532), .A2(n5427), .Y(n5562) );
  NAND3X0_RVT U4855 ( .A1(n5564), .A2(n5565), .A3(n5566), .Y(n4869) );
  NAND2X0_RVT U4856 ( .A1(n5545), .A2(n5431), .Y(n5566) );
  NAND2X0_RVT U4857 ( .A1(n5546), .A2(n5147), .Y(n5565) );
  NAND2X0_RVT U4858 ( .A1(n5567), .A2(n5548), .Y(n5564) );
  NAND3X0_RVT U4859 ( .A1(n5568), .A2(n5569), .A3(n5435), .Y(n5567) );
  NAND2X0_RVT U4860 ( .A1(n5551), .A2(n5436), .Y(n5569) );
  NAND2X0_RVT U4861 ( .A1(n5532), .A2(n5437), .Y(n5568) );
  NAND3X0_RVT U4862 ( .A1(n5570), .A2(n5571), .A3(n5572), .Y(n4868) );
  NAND2X0_RVT U4863 ( .A1(n5545), .A2(n5441), .Y(n5572) );
  NAND2X0_RVT U4864 ( .A1(n5546), .A2(n5152), .Y(n5571) );
  NAND2X0_RVT U4865 ( .A1(n5573), .A2(n5548), .Y(n5570) );
  NAND3X0_RVT U4866 ( .A1(n5574), .A2(n5575), .A3(n5445), .Y(n5573) );
  NAND2X0_RVT U4867 ( .A1(n5551), .A2(n5446), .Y(n5575) );
  NAND2X0_RVT U4868 ( .A1(n5447), .A2(n5532), .Y(n5574) );
  NAND3X0_RVT U4869 ( .A1(n5576), .A2(n5577), .A3(n5578), .Y(n4867) );
  NAND2X0_RVT U4870 ( .A1(n5545), .A2(n5451), .Y(n5578) );
  NAND2X0_RVT U4871 ( .A1(n5546), .A2(n5157), .Y(n5577) );
  NAND2X0_RVT U4872 ( .A1(n5579), .A2(n5548), .Y(n5576) );
  NAND3X0_RVT U4873 ( .A1(n5580), .A2(n5581), .A3(n5455), .Y(n5579) );
  NAND2X0_RVT U4874 ( .A1(n5551), .A2(n5456), .Y(n5581) );
  NAND2X0_RVT U4875 ( .A1(n5532), .A2(n5457), .Y(n5580) );
  NAND3X0_RVT U4876 ( .A1(n5582), .A2(n5583), .A3(n5584), .Y(n4866) );
  NAND2X0_RVT U4877 ( .A1(n5545), .A2(n5461), .Y(n5584) );
  NAND2X0_RVT U4878 ( .A1(n5546), .A2(n5162), .Y(n5583) );
  NAND2X0_RVT U4879 ( .A1(n5585), .A2(n5548), .Y(n5582) );
  NAND3X0_RVT U4880 ( .A1(n5586), .A2(n5587), .A3(n5465), .Y(n5585) );
  NAND2X0_RVT U4881 ( .A1(n5551), .A2(n5466), .Y(n5587) );
  NAND2X0_RVT U4882 ( .A1(n5532), .A2(n5467), .Y(n5586) );
  NAND3X0_RVT U4883 ( .A1(n5588), .A2(n5589), .A3(n5590), .Y(n4865) );
  NAND2X0_RVT U4884 ( .A1(n5545), .A2(n5329), .Y(n5590) );
  AND2X1_RVT U4885 ( .A1(n5480), .A2(n5548), .Y(n5545) );
  NAND2X0_RVT U4886 ( .A1(n5546), .A2(n5168), .Y(n5589) );
  INVX0_RVT U4887 ( .A(n5548), .Y(n5546) );
  NAND2X0_RVT U4888 ( .A1(n5591), .A2(n5548), .Y(n5588) );
  NAND3X0_RVT U4889 ( .A1(n5592), .A2(n5593), .A3(n5594), .Y(n5548) );
  NAND2X0_RVT U4890 ( .A1(n5595), .A2(n5359), .Y(n5594) );
  NAND2X0_RVT U4891 ( .A1(n5476), .A2(n5478), .Y(n5593) );
  NAND2X0_RVT U4892 ( .A1(n5596), .A2(n5479), .Y(n5592) );
  NAND3X0_RVT U4893 ( .A1(n5597), .A2(n5598), .A3(n5334), .Y(n5591) );
  NAND2X0_RVT U4894 ( .A1(n5551), .A2(n5335), .Y(n5598) );
  INVX0_RVT U4895 ( .A(n5478), .Y(n5551) );
  NAND2X0_RVT U4896 ( .A1(n5599), .A2(n5600), .Y(n5478) );
  NAND2X0_RVT U4897 ( .A1(n5338), .A2(n5532), .Y(n5597) );
  NAND3X0_RVT U4898 ( .A1(n5601), .A2(n5602), .A3(n5603), .Y(n4864) );
  NAND2X0_RVT U4899 ( .A1(n5604), .A2(n5397), .Y(n5603) );
  NAND2X0_RVT U4900 ( .A1(n5605), .A2(n5136), .Y(n5602) );
  NAND2X0_RVT U4901 ( .A1(n5606), .A2(n5607), .Y(n5601) );
  NAND3X0_RVT U4902 ( .A1(n5608), .A2(n5609), .A3(n5403), .Y(n5606) );
  NAND2X0_RVT U4903 ( .A1(n5610), .A2(n5404), .Y(n5609) );
  NAND2X0_RVT U4904 ( .A1(n5480), .A2(n5407), .Y(n5608) );
  NAND3X0_RVT U4905 ( .A1(n5611), .A2(n5612), .A3(n5613), .Y(n4863) );
  NAND2X0_RVT U4906 ( .A1(n5604), .A2(n5411), .Y(n5613) );
  NAND2X0_RVT U4907 ( .A1(n5605), .A2(n5141), .Y(n5612) );
  NAND2X0_RVT U4908 ( .A1(n5614), .A2(n5607), .Y(n5611) );
  NAND3X0_RVT U4909 ( .A1(n5615), .A2(n5616), .A3(n5415), .Y(n5614) );
  NAND2X0_RVT U4910 ( .A1(n5610), .A2(n5416), .Y(n5616) );
  NAND2X0_RVT U4911 ( .A1(n5480), .A2(n5417), .Y(n5615) );
  NAND3X0_RVT U4912 ( .A1(n5617), .A2(n5618), .A3(n5619), .Y(n4862) );
  NAND2X0_RVT U4913 ( .A1(n5604), .A2(n5421), .Y(n5619) );
  NAND2X0_RVT U4914 ( .A1(n5605), .A2(n5146), .Y(n5618) );
  NAND2X0_RVT U4915 ( .A1(n5620), .A2(n5607), .Y(n5617) );
  NAND3X0_RVT U4916 ( .A1(n5621), .A2(n5622), .A3(n5425), .Y(n5620) );
  NAND2X0_RVT U4917 ( .A1(n5610), .A2(n5426), .Y(n5622) );
  NAND2X0_RVT U4918 ( .A1(n5480), .A2(n5427), .Y(n5621) );
  NAND3X0_RVT U4919 ( .A1(n5623), .A2(n5624), .A3(n5625), .Y(n4861) );
  NAND2X0_RVT U4920 ( .A1(n5604), .A2(n5431), .Y(n5625) );
  NAND2X0_RVT U4921 ( .A1(n5605), .A2(n5151), .Y(n5624) );
  NAND2X0_RVT U4922 ( .A1(n5626), .A2(n5607), .Y(n5623) );
  NAND3X0_RVT U4923 ( .A1(n5627), .A2(n5628), .A3(n5435), .Y(n5626) );
  NAND2X0_RVT U4924 ( .A1(n5610), .A2(n5436), .Y(n5628) );
  NAND2X0_RVT U4925 ( .A1(n5480), .A2(n5437), .Y(n5627) );
  NAND3X0_RVT U4926 ( .A1(n5629), .A2(n5630), .A3(n5631), .Y(n4860) );
  NAND2X0_RVT U4927 ( .A1(n5604), .A2(n5441), .Y(n5631) );
  NAND2X0_RVT U4928 ( .A1(n5605), .A2(n5156), .Y(n5630) );
  NAND2X0_RVT U4929 ( .A1(n5632), .A2(n5607), .Y(n5629) );
  NAND3X0_RVT U4930 ( .A1(n5633), .A2(n5634), .A3(n5445), .Y(n5632) );
  NAND2X0_RVT U4931 ( .A1(n5610), .A2(n5446), .Y(n5634) );
  NAND2X0_RVT U4932 ( .A1(n5447), .A2(n5480), .Y(n5633) );
  NAND3X0_RVT U4933 ( .A1(n5635), .A2(n5636), .A3(n5637), .Y(n4859) );
  NAND2X0_RVT U4934 ( .A1(n5604), .A2(n5451), .Y(n5637) );
  NAND2X0_RVT U4935 ( .A1(n5605), .A2(n5161), .Y(n5636) );
  NAND2X0_RVT U4936 ( .A1(n5638), .A2(n5607), .Y(n5635) );
  NAND3X0_RVT U4937 ( .A1(n5639), .A2(n5640), .A3(n5455), .Y(n5638) );
  NAND2X0_RVT U4938 ( .A1(n5610), .A2(n5456), .Y(n5640) );
  NAND2X0_RVT U4939 ( .A1(n5480), .A2(n5457), .Y(n5639) );
  NAND3X0_RVT U4940 ( .A1(n5641), .A2(n5642), .A3(n5643), .Y(n4858) );
  NAND2X0_RVT U4941 ( .A1(n5604), .A2(n5461), .Y(n5643) );
  NAND2X0_RVT U4942 ( .A1(n5605), .A2(n5166), .Y(n5642) );
  NAND2X0_RVT U4943 ( .A1(n5644), .A2(n5607), .Y(n5641) );
  NAND3X0_RVT U4944 ( .A1(n5645), .A2(n5646), .A3(n5465), .Y(n5644) );
  NAND2X0_RVT U4945 ( .A1(n5610), .A2(n5466), .Y(n5646) );
  NAND2X0_RVT U4946 ( .A1(n5480), .A2(n5467), .Y(n5645) );
  NAND3X0_RVT U4947 ( .A1(n5647), .A2(n5648), .A3(n5649), .Y(n4857) );
  NAND2X0_RVT U4948 ( .A1(n5604), .A2(n5329), .Y(n5649) );
  AND2X1_RVT U4949 ( .A1(n5539), .A2(n5607), .Y(n5604) );
  NAND2X0_RVT U4950 ( .A1(n5605), .A2(n5172), .Y(n5648) );
  INVX0_RVT U4951 ( .A(n5607), .Y(n5605) );
  NAND2X0_RVT U4952 ( .A1(n5650), .A2(n5607), .Y(n5647) );
  NAND3X0_RVT U4953 ( .A1(n5651), .A2(n5652), .A3(n5653), .Y(n5607) );
  NAND2X0_RVT U4954 ( .A1(n5654), .A2(n5359), .Y(n5653) );
  NAND2X0_RVT U4955 ( .A1(n5476), .A2(n5538), .Y(n5652) );
  NAND2X0_RVT U4956 ( .A1(n5655), .A2(n5479), .Y(n5651) );
  NAND3X0_RVT U4957 ( .A1(n5656), .A2(n5657), .A3(n5334), .Y(n5650) );
  NAND2X0_RVT U4958 ( .A1(n5610), .A2(n5335), .Y(n5657) );
  INVX0_RVT U4959 ( .A(n5538), .Y(n5610) );
  NAND2X0_RVT U4960 ( .A1(n5658), .A2(n5600), .Y(n5538) );
  NAND2X0_RVT U4961 ( .A1(n5480), .A2(n5338), .Y(n5656) );
  INVX0_RVT U4962 ( .A(n5600), .Y(n5480) );
  NAND2X0_RVT U4963 ( .A1(n5659), .A2(n5660), .Y(n5600) );
  NAND3X0_RVT U4964 ( .A1(n5661), .A2(n5662), .A3(n5663), .Y(n4856) );
  NAND2X0_RVT U4965 ( .A1(n5664), .A2(n5397), .Y(n5663) );
  NAND2X0_RVT U4966 ( .A1(n5665), .A2(n5134), .Y(n5662) );
  NAND2X0_RVT U4967 ( .A1(n5666), .A2(n5667), .Y(n5661) );
  NAND3X0_RVT U4968 ( .A1(n5668), .A2(n5669), .A3(n5403), .Y(n5666) );
  NAND2X0_RVT U4969 ( .A1(n5670), .A2(n5404), .Y(n5669) );
  NAND2X0_RVT U4970 ( .A1(n5539), .A2(n5407), .Y(n5668) );
  NAND3X0_RVT U4971 ( .A1(n5671), .A2(n5672), .A3(n5673), .Y(n4855) );
  NAND2X0_RVT U4972 ( .A1(n5664), .A2(n5411), .Y(n5673) );
  NAND2X0_RVT U4973 ( .A1(n5665), .A2(n5139), .Y(n5672) );
  NAND2X0_RVT U4974 ( .A1(n5674), .A2(n5667), .Y(n5671) );
  NAND3X0_RVT U4975 ( .A1(n5675), .A2(n5676), .A3(n5415), .Y(n5674) );
  NAND2X0_RVT U4976 ( .A1(n5670), .A2(n5416), .Y(n5676) );
  NAND2X0_RVT U4977 ( .A1(n5539), .A2(n5417), .Y(n5675) );
  NAND3X0_RVT U4978 ( .A1(n5677), .A2(n5678), .A3(n5679), .Y(n4854) );
  NAND2X0_RVT U4979 ( .A1(n5664), .A2(n5421), .Y(n5679) );
  NAND2X0_RVT U4980 ( .A1(n5665), .A2(n5144), .Y(n5678) );
  NAND2X0_RVT U4981 ( .A1(n5680), .A2(n5667), .Y(n5677) );
  NAND3X0_RVT U4982 ( .A1(n5681), .A2(n5682), .A3(n5425), .Y(n5680) );
  NAND2X0_RVT U4983 ( .A1(n5670), .A2(n5426), .Y(n5682) );
  NAND2X0_RVT U4984 ( .A1(n5539), .A2(n5427), .Y(n5681) );
  NAND3X0_RVT U4985 ( .A1(n5683), .A2(n5684), .A3(n5685), .Y(n4853) );
  NAND2X0_RVT U4986 ( .A1(n5664), .A2(n5431), .Y(n5685) );
  NAND2X0_RVT U4987 ( .A1(n5665), .A2(n5149), .Y(n5684) );
  NAND2X0_RVT U4988 ( .A1(n5686), .A2(n5667), .Y(n5683) );
  NAND3X0_RVT U4989 ( .A1(n5687), .A2(n5688), .A3(n5435), .Y(n5686) );
  NAND2X0_RVT U4990 ( .A1(n5670), .A2(n5436), .Y(n5688) );
  NAND2X0_RVT U4991 ( .A1(n5539), .A2(n5437), .Y(n5687) );
  NAND3X0_RVT U4992 ( .A1(n5689), .A2(n5690), .A3(n5691), .Y(n4852) );
  NAND2X0_RVT U4993 ( .A1(n5664), .A2(n5441), .Y(n5691) );
  NAND2X0_RVT U4994 ( .A1(n5665), .A2(n5154), .Y(n5690) );
  NAND2X0_RVT U4995 ( .A1(n5692), .A2(n5667), .Y(n5689) );
  NAND3X0_RVT U4996 ( .A1(n5693), .A2(n5694), .A3(n5445), .Y(n5692) );
  NAND2X0_RVT U4997 ( .A1(n5670), .A2(n5446), .Y(n5694) );
  NAND2X0_RVT U4998 ( .A1(n5539), .A2(n5447), .Y(n5693) );
  NAND3X0_RVT U4999 ( .A1(n5695), .A2(n5696), .A3(n5697), .Y(n4851) );
  NAND2X0_RVT U5000 ( .A1(n5664), .A2(n5451), .Y(n5697) );
  NAND2X0_RVT U5001 ( .A1(n5665), .A2(n5159), .Y(n5696) );
  NAND2X0_RVT U5002 ( .A1(n5698), .A2(n5667), .Y(n5695) );
  NAND3X0_RVT U5003 ( .A1(n5699), .A2(n5700), .A3(n5455), .Y(n5698) );
  NAND2X0_RVT U5004 ( .A1(n5670), .A2(n5456), .Y(n5700) );
  NAND2X0_RVT U5005 ( .A1(n5539), .A2(n5457), .Y(n5699) );
  NAND3X0_RVT U5006 ( .A1(n5701), .A2(n5702), .A3(n5703), .Y(n4850) );
  NAND2X0_RVT U5007 ( .A1(n5664), .A2(n5461), .Y(n5703) );
  NAND2X0_RVT U5008 ( .A1(n5665), .A2(n5164), .Y(n5702) );
  NAND2X0_RVT U5009 ( .A1(n5704), .A2(n5667), .Y(n5701) );
  NAND3X0_RVT U5010 ( .A1(n5705), .A2(n5706), .A3(n5465), .Y(n5704) );
  NAND2X0_RVT U5011 ( .A1(n5670), .A2(n5466), .Y(n5706) );
  NAND2X0_RVT U5012 ( .A1(n5539), .A2(n5467), .Y(n5705) );
  NAND3X0_RVT U5013 ( .A1(n5707), .A2(n5708), .A3(n5709), .Y(n4849) );
  NAND2X0_RVT U5014 ( .A1(n5664), .A2(n5329), .Y(n5709) );
  AND2X1_RVT U5015 ( .A1(n5595), .A2(n5667), .Y(n5664) );
  NAND2X0_RVT U5016 ( .A1(n5665), .A2(n5169), .Y(n5708) );
  INVX0_RVT U5017 ( .A(n5667), .Y(n5665) );
  NAND2X0_RVT U5018 ( .A1(n5710), .A2(n5667), .Y(n5707) );
  NAND3X0_RVT U5019 ( .A1(n5711), .A2(n5712), .A3(n5713), .Y(n5667) );
  NAND2X0_RVT U5020 ( .A1(n5714), .A2(n5359), .Y(n5713) );
  NAND2X0_RVT U5021 ( .A1(n5476), .A2(n5596), .Y(n5712) );
  NAND2X0_RVT U5022 ( .A1(n5715), .A2(n5479), .Y(n5711) );
  NAND3X0_RVT U5023 ( .A1(n5716), .A2(n5717), .A3(n5334), .Y(n5710) );
  NAND2X0_RVT U5024 ( .A1(n5670), .A2(n5335), .Y(n5717) );
  INVX0_RVT U5025 ( .A(n5596), .Y(n5670) );
  NAND2X0_RVT U5026 ( .A1(n5718), .A2(n5658), .Y(n5596) );
  NAND2X0_RVT U5027 ( .A1(n5539), .A2(n5338), .Y(n5716) );
  INVX0_RVT U5028 ( .A(n5658), .Y(n5539) );
  NAND2X0_RVT U5029 ( .A1(n5719), .A2(n5660), .Y(n5658) );
  NAND3X0_RVT U5030 ( .A1(n5720), .A2(n5721), .A3(n5722), .Y(n4848) );
  NAND2X0_RVT U5031 ( .A1(n5723), .A2(n5397), .Y(n5722) );
  NAND2X0_RVT U5032 ( .A1(n5724), .A2(n4997), .Y(n5721) );
  NAND2X0_RVT U5033 ( .A1(n5725), .A2(n5726), .Y(n5720) );
  NAND3X0_RVT U5034 ( .A1(n5727), .A2(n5728), .A3(n5403), .Y(n5725) );
  NAND2X0_RVT U5035 ( .A1(n5729), .A2(n5404), .Y(n5728) );
  NAND2X0_RVT U5036 ( .A1(n5595), .A2(n5407), .Y(n5727) );
  NAND3X0_RVT U5037 ( .A1(n5730), .A2(n5731), .A3(n5732), .Y(n4847) );
  NAND2X0_RVT U5038 ( .A1(n5723), .A2(n5411), .Y(n5732) );
  NAND2X0_RVT U5039 ( .A1(n5724), .A2(n5004), .Y(n5731) );
  NAND2X0_RVT U5040 ( .A1(n5733), .A2(n5726), .Y(n5730) );
  NAND3X0_RVT U5041 ( .A1(n5734), .A2(n5735), .A3(n5415), .Y(n5733) );
  NAND2X0_RVT U5042 ( .A1(n5729), .A2(n5416), .Y(n5735) );
  NAND2X0_RVT U5043 ( .A1(n5595), .A2(n5417), .Y(n5734) );
  NAND3X0_RVT U5044 ( .A1(n5736), .A2(n5737), .A3(n5738), .Y(n4846) );
  NAND2X0_RVT U5045 ( .A1(n5723), .A2(n5421), .Y(n5738) );
  NAND2X0_RVT U5046 ( .A1(n5724), .A2(n5011), .Y(n5737) );
  NAND2X0_RVT U5047 ( .A1(n5739), .A2(n5726), .Y(n5736) );
  NAND3X0_RVT U5048 ( .A1(n5740), .A2(n5741), .A3(n5425), .Y(n5739) );
  NAND2X0_RVT U5049 ( .A1(n5729), .A2(n5426), .Y(n5741) );
  NAND2X0_RVT U5050 ( .A1(n5595), .A2(n5427), .Y(n5740) );
  NAND3X0_RVT U5051 ( .A1(n5742), .A2(n5743), .A3(n5744), .Y(n4845) );
  NAND2X0_RVT U5052 ( .A1(n5723), .A2(n5431), .Y(n5744) );
  NAND2X0_RVT U5053 ( .A1(n5724), .A2(n5017), .Y(n5743) );
  NAND2X0_RVT U5054 ( .A1(n5745), .A2(n5726), .Y(n5742) );
  NAND3X0_RVT U5055 ( .A1(n5746), .A2(n5747), .A3(n5435), .Y(n5745) );
  NAND2X0_RVT U5056 ( .A1(n5729), .A2(n5436), .Y(n5747) );
  NAND2X0_RVT U5057 ( .A1(n5595), .A2(n5437), .Y(n5746) );
  NAND3X0_RVT U5058 ( .A1(n5748), .A2(n5749), .A3(n5750), .Y(n4844) );
  NAND2X0_RVT U5059 ( .A1(n5723), .A2(n5441), .Y(n5750) );
  NAND2X0_RVT U5060 ( .A1(n5724), .A2(n5024), .Y(n5749) );
  NAND2X0_RVT U5061 ( .A1(n5751), .A2(n5726), .Y(n5748) );
  NAND3X0_RVT U5062 ( .A1(n5752), .A2(n5753), .A3(n5445), .Y(n5751) );
  NAND2X0_RVT U5063 ( .A1(n5729), .A2(n5446), .Y(n5753) );
  NAND2X0_RVT U5064 ( .A1(n5595), .A2(n5447), .Y(n5752) );
  NAND3X0_RVT U5065 ( .A1(n5754), .A2(n5755), .A3(n5756), .Y(n4843) );
  NAND2X0_RVT U5066 ( .A1(n5723), .A2(n5451), .Y(n5756) );
  NAND2X0_RVT U5067 ( .A1(n5724), .A2(n5031), .Y(n5755) );
  NAND2X0_RVT U5068 ( .A1(n5757), .A2(n5726), .Y(n5754) );
  NAND3X0_RVT U5069 ( .A1(n5758), .A2(n5759), .A3(n5455), .Y(n5757) );
  NAND2X0_RVT U5070 ( .A1(n5729), .A2(n5456), .Y(n5759) );
  NAND2X0_RVT U5071 ( .A1(n5595), .A2(n5457), .Y(n5758) );
  NAND3X0_RVT U5072 ( .A1(n5760), .A2(n5761), .A3(n5762), .Y(n4842) );
  NAND2X0_RVT U5073 ( .A1(n5723), .A2(n5461), .Y(n5762) );
  NAND2X0_RVT U5074 ( .A1(n5724), .A2(n5038), .Y(n5761) );
  NAND2X0_RVT U5075 ( .A1(n5763), .A2(n5726), .Y(n5760) );
  NAND3X0_RVT U5076 ( .A1(n5764), .A2(n5765), .A3(n5465), .Y(n5763) );
  NAND2X0_RVT U5077 ( .A1(n5729), .A2(n5466), .Y(n5765) );
  NAND2X0_RVT U5078 ( .A1(n5595), .A2(n5467), .Y(n5764) );
  NAND3X0_RVT U5079 ( .A1(n5766), .A2(n5767), .A3(n5768), .Y(n4841) );
  NAND2X0_RVT U5080 ( .A1(n5723), .A2(n5329), .Y(n5768) );
  AND2X1_RVT U5081 ( .A1(n5654), .A2(n5726), .Y(n5723) );
  NAND2X0_RVT U5082 ( .A1(n5724), .A2(n5043), .Y(n5767) );
  INVX0_RVT U5083 ( .A(n5726), .Y(n5724) );
  NAND2X0_RVT U5084 ( .A1(n5769), .A2(n5726), .Y(n5766) );
  NAND3X0_RVT U5085 ( .A1(n5770), .A2(n5771), .A3(n5772), .Y(n5726) );
  NAND2X0_RVT U5086 ( .A1(n5773), .A2(n5359), .Y(n5772) );
  NAND2X0_RVT U5087 ( .A1(n5476), .A2(n5655), .Y(n5771) );
  NAND2X0_RVT U5088 ( .A1(n5774), .A2(n5479), .Y(n5770) );
  NAND3X0_RVT U5089 ( .A1(n5775), .A2(n5776), .A3(n5334), .Y(n5769) );
  NAND2X0_RVT U5090 ( .A1(n5729), .A2(n5335), .Y(n5776) );
  INVX0_RVT U5091 ( .A(n5655), .Y(n5729) );
  NAND2X0_RVT U5092 ( .A1(n5777), .A2(n5718), .Y(n5655) );
  NAND2X0_RVT U5093 ( .A1(n5595), .A2(n5338), .Y(n5775) );
  INVX0_RVT U5094 ( .A(n5718), .Y(n5595) );
  NAND2X0_RVT U5095 ( .A1(n5778), .A2(n5659), .Y(n5718) );
  NAND3X0_RVT U5096 ( .A1(n5779), .A2(n5780), .A3(n5781), .Y(n4840) );
  NAND2X0_RVT U5097 ( .A1(n5782), .A2(n5397), .Y(n5781) );
  NAND2X0_RVT U5098 ( .A1(n5783), .A2(n5000), .Y(n5780) );
  NAND2X0_RVT U5099 ( .A1(n5784), .A2(n5785), .Y(n5779) );
  NAND3X0_RVT U5100 ( .A1(n5786), .A2(n5787), .A3(n5403), .Y(n5784) );
  NAND2X0_RVT U5101 ( .A1(n5788), .A2(n5404), .Y(n5787) );
  NAND2X0_RVT U5102 ( .A1(n5654), .A2(n5407), .Y(n5786) );
  NAND3X0_RVT U5103 ( .A1(n5789), .A2(n5790), .A3(n5791), .Y(n4839) );
  NAND2X0_RVT U5104 ( .A1(n5782), .A2(n5411), .Y(n5791) );
  NAND2X0_RVT U5105 ( .A1(n5783), .A2(n5007), .Y(n5790) );
  NAND2X0_RVT U5106 ( .A1(n5792), .A2(n5785), .Y(n5789) );
  NAND3X0_RVT U5107 ( .A1(n5793), .A2(n5794), .A3(n5415), .Y(n5792) );
  NAND2X0_RVT U5108 ( .A1(n5788), .A2(n5416), .Y(n5794) );
  NAND2X0_RVT U5109 ( .A1(n5654), .A2(n5417), .Y(n5793) );
  NAND3X0_RVT U5110 ( .A1(n5795), .A2(n5796), .A3(n5797), .Y(n4838) );
  NAND2X0_RVT U5111 ( .A1(n5782), .A2(n5421), .Y(n5797) );
  NAND2X0_RVT U5112 ( .A1(n5783), .A2(n5014), .Y(n5796) );
  NAND2X0_RVT U5113 ( .A1(n5798), .A2(n5785), .Y(n5795) );
  NAND3X0_RVT U5114 ( .A1(n5799), .A2(n5800), .A3(n5425), .Y(n5798) );
  NAND2X0_RVT U5115 ( .A1(n5788), .A2(n5426), .Y(n5800) );
  NAND2X0_RVT U5116 ( .A1(n5654), .A2(n5427), .Y(n5799) );
  NAND3X0_RVT U5117 ( .A1(n5801), .A2(n5802), .A3(n5803), .Y(n4837) );
  NAND2X0_RVT U5118 ( .A1(n5782), .A2(n5431), .Y(n5803) );
  NAND2X0_RVT U5119 ( .A1(n5783), .A2(n5020), .Y(n5802) );
  NAND2X0_RVT U5120 ( .A1(n5804), .A2(n5785), .Y(n5801) );
  NAND3X0_RVT U5121 ( .A1(n5805), .A2(n5806), .A3(n5435), .Y(n5804) );
  NAND2X0_RVT U5122 ( .A1(n5788), .A2(n5436), .Y(n5806) );
  NAND2X0_RVT U5123 ( .A1(n5654), .A2(n5437), .Y(n5805) );
  NAND3X0_RVT U5124 ( .A1(n5807), .A2(n5808), .A3(n5809), .Y(n4836) );
  NAND2X0_RVT U5125 ( .A1(n5782), .A2(n5441), .Y(n5809) );
  NAND2X0_RVT U5126 ( .A1(n5783), .A2(n5027), .Y(n5808) );
  NAND2X0_RVT U5127 ( .A1(n5810), .A2(n5785), .Y(n5807) );
  NAND3X0_RVT U5128 ( .A1(n5811), .A2(n5812), .A3(n5445), .Y(n5810) );
  NAND2X0_RVT U5129 ( .A1(n5788), .A2(n5446), .Y(n5812) );
  NAND2X0_RVT U5130 ( .A1(n5654), .A2(n5447), .Y(n5811) );
  NAND3X0_RVT U5131 ( .A1(n5813), .A2(n5814), .A3(n5815), .Y(n4835) );
  NAND2X0_RVT U5132 ( .A1(n5782), .A2(n5451), .Y(n5815) );
  NAND2X0_RVT U5133 ( .A1(n5783), .A2(n5034), .Y(n5814) );
  NAND2X0_RVT U5134 ( .A1(n5816), .A2(n5785), .Y(n5813) );
  NAND3X0_RVT U5135 ( .A1(n5817), .A2(n5818), .A3(n5455), .Y(n5816) );
  NAND2X0_RVT U5136 ( .A1(n5788), .A2(n5456), .Y(n5818) );
  NAND2X0_RVT U5137 ( .A1(n5654), .A2(n5457), .Y(n5817) );
  NAND3X0_RVT U5138 ( .A1(n5819), .A2(n5820), .A3(n5821), .Y(n4834) );
  NAND2X0_RVT U5139 ( .A1(n5782), .A2(n5461), .Y(n5821) );
  NAND2X0_RVT U5140 ( .A1(n5783), .A2(n5041), .Y(n5820) );
  NAND2X0_RVT U5141 ( .A1(n5822), .A2(n5785), .Y(n5819) );
  NAND3X0_RVT U5142 ( .A1(n5823), .A2(n5824), .A3(n5465), .Y(n5822) );
  NAND2X0_RVT U5143 ( .A1(n5788), .A2(n5466), .Y(n5824) );
  NAND2X0_RVT U5144 ( .A1(n5654), .A2(n5467), .Y(n5823) );
  NAND3X0_RVT U5145 ( .A1(n5825), .A2(n5826), .A3(n5827), .Y(n4833) );
  NAND2X0_RVT U5146 ( .A1(n5782), .A2(n5329), .Y(n5827) );
  AND2X1_RVT U5147 ( .A1(n5714), .A2(n5785), .Y(n5782) );
  NAND2X0_RVT U5148 ( .A1(n5783), .A2(n5046), .Y(n5826) );
  INVX0_RVT U5149 ( .A(n5785), .Y(n5783) );
  NAND2X0_RVT U5150 ( .A1(n5828), .A2(n5785), .Y(n5825) );
  NAND3X0_RVT U5151 ( .A1(n5829), .A2(n5830), .A3(n5831), .Y(n5785) );
  NAND2X0_RVT U5152 ( .A1(n5832), .A2(n5359), .Y(n5831) );
  NAND2X0_RVT U5153 ( .A1(n5476), .A2(n5715), .Y(n5830) );
  NAND2X0_RVT U5154 ( .A1(n5833), .A2(n5479), .Y(n5829) );
  NAND3X0_RVT U5155 ( .A1(n5834), .A2(n5835), .A3(n5334), .Y(n5828) );
  NAND2X0_RVT U5156 ( .A1(n5788), .A2(n5335), .Y(n5835) );
  INVX0_RVT U5157 ( .A(n5715), .Y(n5788) );
  NAND2X0_RVT U5158 ( .A1(n5836), .A2(n5777), .Y(n5715) );
  NAND2X0_RVT U5159 ( .A1(n5654), .A2(n5338), .Y(n5834) );
  INVX0_RVT U5160 ( .A(n5777), .Y(n5654) );
  NAND2X0_RVT U5161 ( .A1(n5778), .A2(n5719), .Y(n5777) );
  NAND3X0_RVT U5162 ( .A1(n5837), .A2(n5838), .A3(n5839), .Y(n4832) );
  NAND2X0_RVT U5163 ( .A1(n5840), .A2(n5397), .Y(n5839) );
  NAND2X0_RVT U5164 ( .A1(n5841), .A2(n5002), .Y(n5838) );
  NAND2X0_RVT U5165 ( .A1(n5842), .A2(n5843), .Y(n5837) );
  NAND3X0_RVT U5166 ( .A1(n5844), .A2(n5845), .A3(n5403), .Y(n5842) );
  NAND2X0_RVT U5167 ( .A1(n5846), .A2(n5404), .Y(n5845) );
  NAND2X0_RVT U5168 ( .A1(n5714), .A2(n5407), .Y(n5844) );
  NAND3X0_RVT U5169 ( .A1(n5847), .A2(n5848), .A3(n5849), .Y(n4831) );
  NAND2X0_RVT U5170 ( .A1(n5840), .A2(n5411), .Y(n5849) );
  NAND2X0_RVT U5171 ( .A1(n5841), .A2(n5009), .Y(n5848) );
  NAND2X0_RVT U5172 ( .A1(n5850), .A2(n5843), .Y(n5847) );
  NAND3X0_RVT U5173 ( .A1(n5851), .A2(n5852), .A3(n5415), .Y(n5850) );
  NAND2X0_RVT U5174 ( .A1(n5846), .A2(n5416), .Y(n5852) );
  NAND2X0_RVT U5175 ( .A1(n5714), .A2(n5417), .Y(n5851) );
  NAND3X0_RVT U5176 ( .A1(n5853), .A2(n5854), .A3(n5855), .Y(n4830) );
  NAND2X0_RVT U5177 ( .A1(n5840), .A2(n5421), .Y(n5855) );
  NAND2X0_RVT U5178 ( .A1(n5841), .A2(n5108), .Y(n5854) );
  NAND2X0_RVT U5179 ( .A1(n5856), .A2(n5843), .Y(n5853) );
  NAND3X0_RVT U5180 ( .A1(n5857), .A2(n5858), .A3(n5425), .Y(n5856) );
  NAND2X0_RVT U5181 ( .A1(n5846), .A2(n5426), .Y(n5858) );
  NAND2X0_RVT U5182 ( .A1(n5714), .A2(n5427), .Y(n5857) );
  NAND3X0_RVT U5183 ( .A1(n5859), .A2(n5860), .A3(n5861), .Y(n4829) );
  NAND2X0_RVT U5184 ( .A1(n5840), .A2(n5431), .Y(n5861) );
  NAND2X0_RVT U5185 ( .A1(n5841), .A2(n5022), .Y(n5860) );
  NAND2X0_RVT U5186 ( .A1(n5862), .A2(n5843), .Y(n5859) );
  NAND3X0_RVT U5187 ( .A1(n5863), .A2(n5864), .A3(n5435), .Y(n5862) );
  NAND2X0_RVT U5188 ( .A1(n5846), .A2(n5436), .Y(n5864) );
  NAND2X0_RVT U5189 ( .A1(n5714), .A2(n5437), .Y(n5863) );
  NAND3X0_RVT U5190 ( .A1(n5865), .A2(n5866), .A3(n5867), .Y(n4828) );
  NAND2X0_RVT U5191 ( .A1(n5840), .A2(n5441), .Y(n5867) );
  NAND2X0_RVT U5192 ( .A1(n5841), .A2(n5029), .Y(n5866) );
  NAND2X0_RVT U5193 ( .A1(n5868), .A2(n5843), .Y(n5865) );
  NAND3X0_RVT U5194 ( .A1(n5869), .A2(n5870), .A3(n5445), .Y(n5868) );
  NAND2X0_RVT U5195 ( .A1(n5846), .A2(n5446), .Y(n5870) );
  NAND2X0_RVT U5196 ( .A1(n5714), .A2(n5447), .Y(n5869) );
  NAND3X0_RVT U5197 ( .A1(n5871), .A2(n5872), .A3(n5873), .Y(n4827) );
  NAND2X0_RVT U5198 ( .A1(n5840), .A2(n5451), .Y(n5873) );
  NAND2X0_RVT U5199 ( .A1(n5841), .A2(n5036), .Y(n5872) );
  NAND2X0_RVT U5200 ( .A1(n5874), .A2(n5843), .Y(n5871) );
  NAND3X0_RVT U5201 ( .A1(n5875), .A2(n5876), .A3(n5455), .Y(n5874) );
  NAND2X0_RVT U5202 ( .A1(n5846), .A2(n5456), .Y(n5876) );
  NAND2X0_RVT U5203 ( .A1(n5714), .A2(n5457), .Y(n5875) );
  NAND3X0_RVT U5204 ( .A1(n5877), .A2(n5878), .A3(n5879), .Y(n4826) );
  NAND2X0_RVT U5205 ( .A1(n5840), .A2(n5461), .Y(n5879) );
  NAND2X0_RVT U5206 ( .A1(n5841), .A2(n5109), .Y(n5878) );
  NAND2X0_RVT U5207 ( .A1(n5880), .A2(n5843), .Y(n5877) );
  NAND3X0_RVT U5208 ( .A1(n5881), .A2(n5882), .A3(n5465), .Y(n5880) );
  NAND2X0_RVT U5209 ( .A1(n5846), .A2(n5466), .Y(n5882) );
  NAND2X0_RVT U5210 ( .A1(n5714), .A2(n5467), .Y(n5881) );
  NAND3X0_RVT U5211 ( .A1(n5883), .A2(n5884), .A3(n5885), .Y(n4825) );
  NAND2X0_RVT U5212 ( .A1(n5840), .A2(n5329), .Y(n5885) );
  AND2X1_RVT U5213 ( .A1(n5773), .A2(n5843), .Y(n5840) );
  NAND2X0_RVT U5214 ( .A1(n5841), .A2(n5050), .Y(n5884) );
  INVX0_RVT U5215 ( .A(n5843), .Y(n5841) );
  NAND2X0_RVT U5216 ( .A1(n5886), .A2(n5843), .Y(n5883) );
  NAND3X0_RVT U5217 ( .A1(n5887), .A2(n5888), .A3(n5889), .Y(n5843) );
  NAND2X0_RVT U5218 ( .A1(n5890), .A2(n5359), .Y(n5889) );
  NAND2X0_RVT U5219 ( .A1(n5476), .A2(n5774), .Y(n5888) );
  NAND2X0_RVT U5220 ( .A1(n5891), .A2(n5479), .Y(n5887) );
  NAND3X0_RVT U5221 ( .A1(n5892), .A2(n5893), .A3(n5334), .Y(n5886) );
  NAND2X0_RVT U5222 ( .A1(n5846), .A2(n5335), .Y(n5893) );
  INVX0_RVT U5223 ( .A(n5774), .Y(n5846) );
  NAND2X0_RVT U5224 ( .A1(n5894), .A2(n5836), .Y(n5774) );
  NAND2X0_RVT U5225 ( .A1(n5714), .A2(n5338), .Y(n5892) );
  INVX0_RVT U5226 ( .A(n5836), .Y(n5714) );
  NAND2X0_RVT U5227 ( .A1(n5660), .A2(n5895), .Y(n5836) );
  NAND3X0_RVT U5228 ( .A1(n5896), .A2(n5897), .A3(n5898), .Y(n4824) );
  NAND2X0_RVT U5229 ( .A1(n5899), .A2(n5397), .Y(n5898) );
  NAND2X0_RVT U5230 ( .A1(n5900), .A2(n5135), .Y(n5897) );
  NAND2X0_RVT U5231 ( .A1(n5901), .A2(n5902), .Y(n5896) );
  NAND3X0_RVT U5232 ( .A1(n5903), .A2(n5904), .A3(n5403), .Y(n5901) );
  NAND2X0_RVT U5233 ( .A1(n5905), .A2(n5404), .Y(n5904) );
  NAND2X0_RVT U5234 ( .A1(n5773), .A2(n5407), .Y(n5903) );
  NAND3X0_RVT U5235 ( .A1(n5906), .A2(n5907), .A3(n5908), .Y(n4823) );
  NAND2X0_RVT U5236 ( .A1(n5899), .A2(n5411), .Y(n5908) );
  NAND2X0_RVT U5237 ( .A1(n5900), .A2(n5140), .Y(n5907) );
  NAND2X0_RVT U5238 ( .A1(n5909), .A2(n5902), .Y(n5906) );
  NAND3X0_RVT U5239 ( .A1(n5910), .A2(n5911), .A3(n5415), .Y(n5909) );
  NAND2X0_RVT U5240 ( .A1(n5905), .A2(n5416), .Y(n5911) );
  NAND2X0_RVT U5241 ( .A1(n5773), .A2(n5417), .Y(n5910) );
  NAND3X0_RVT U5242 ( .A1(n5912), .A2(n5913), .A3(n5914), .Y(n4822) );
  NAND2X0_RVT U5243 ( .A1(n5899), .A2(n5421), .Y(n5914) );
  NAND2X0_RVT U5244 ( .A1(n5900), .A2(n5145), .Y(n5913) );
  NAND2X0_RVT U5245 ( .A1(n5915), .A2(n5902), .Y(n5912) );
  NAND3X0_RVT U5246 ( .A1(n5916), .A2(n5917), .A3(n5425), .Y(n5915) );
  NAND2X0_RVT U5247 ( .A1(n5905), .A2(n5426), .Y(n5917) );
  NAND2X0_RVT U5248 ( .A1(n5773), .A2(n5427), .Y(n5916) );
  NAND3X0_RVT U5249 ( .A1(n5918), .A2(n5919), .A3(n5920), .Y(n4821) );
  NAND2X0_RVT U5250 ( .A1(n5899), .A2(n5431), .Y(n5920) );
  NAND2X0_RVT U5251 ( .A1(n5900), .A2(n5150), .Y(n5919) );
  NAND2X0_RVT U5252 ( .A1(n5921), .A2(n5902), .Y(n5918) );
  NAND3X0_RVT U5253 ( .A1(n5922), .A2(n5923), .A3(n5435), .Y(n5921) );
  NAND2X0_RVT U5254 ( .A1(n5905), .A2(n5436), .Y(n5923) );
  NAND2X0_RVT U5255 ( .A1(n5773), .A2(n5437), .Y(n5922) );
  NAND3X0_RVT U5256 ( .A1(n5924), .A2(n5925), .A3(n5926), .Y(n4820) );
  NAND2X0_RVT U5257 ( .A1(n5899), .A2(n5441), .Y(n5926) );
  NAND2X0_RVT U5258 ( .A1(n5900), .A2(n5155), .Y(n5925) );
  NAND2X0_RVT U5259 ( .A1(n5927), .A2(n5902), .Y(n5924) );
  NAND3X0_RVT U5260 ( .A1(n5928), .A2(n5929), .A3(n5445), .Y(n5927) );
  NAND2X0_RVT U5261 ( .A1(n5905), .A2(n5446), .Y(n5929) );
  NAND2X0_RVT U5262 ( .A1(n5773), .A2(n5447), .Y(n5928) );
  NAND3X0_RVT U5263 ( .A1(n5930), .A2(n5931), .A3(n5932), .Y(n4819) );
  NAND2X0_RVT U5264 ( .A1(n5899), .A2(n5451), .Y(n5932) );
  NAND2X0_RVT U5265 ( .A1(n5900), .A2(n5160), .Y(n5931) );
  NAND2X0_RVT U5266 ( .A1(n5933), .A2(n5902), .Y(n5930) );
  NAND3X0_RVT U5267 ( .A1(n5934), .A2(n5935), .A3(n5455), .Y(n5933) );
  NAND2X0_RVT U5268 ( .A1(n5905), .A2(n5456), .Y(n5935) );
  NAND2X0_RVT U5269 ( .A1(n5773), .A2(n5457), .Y(n5934) );
  NAND3X0_RVT U5270 ( .A1(n5936), .A2(n5937), .A3(n5938), .Y(n4818) );
  NAND2X0_RVT U5271 ( .A1(n5899), .A2(n5461), .Y(n5938) );
  NAND2X0_RVT U5272 ( .A1(n5900), .A2(n5165), .Y(n5937) );
  NAND2X0_RVT U5273 ( .A1(n5939), .A2(n5902), .Y(n5936) );
  NAND3X0_RVT U5274 ( .A1(n5940), .A2(n5941), .A3(n5465), .Y(n5939) );
  NAND2X0_RVT U5275 ( .A1(n5905), .A2(n5466), .Y(n5941) );
  NAND2X0_RVT U5276 ( .A1(n5773), .A2(n5467), .Y(n5940) );
  NAND3X0_RVT U5277 ( .A1(n5942), .A2(n5943), .A3(n5944), .Y(n4817) );
  NAND2X0_RVT U5278 ( .A1(n5899), .A2(n5329), .Y(n5944) );
  AND2X1_RVT U5279 ( .A1(n5832), .A2(n5902), .Y(n5899) );
  NAND2X0_RVT U5280 ( .A1(n5900), .A2(n5170), .Y(n5943) );
  INVX0_RVT U5281 ( .A(n5902), .Y(n5900) );
  NAND2X0_RVT U5282 ( .A1(n5945), .A2(n5902), .Y(n5942) );
  NAND3X0_RVT U5283 ( .A1(n5946), .A2(n5947), .A3(n5948), .Y(n5902) );
  NAND2X0_RVT U5284 ( .A1(n5949), .A2(n5359), .Y(n5948) );
  NAND2X0_RVT U5285 ( .A1(n5476), .A2(n5833), .Y(n5947) );
  NAND2X0_RVT U5286 ( .A1(n5950), .A2(n5479), .Y(n5946) );
  NAND3X0_RVT U5287 ( .A1(n5951), .A2(n5952), .A3(n5334), .Y(n5945) );
  NAND2X0_RVT U5288 ( .A1(n5905), .A2(n5335), .Y(n5952) );
  INVX0_RVT U5289 ( .A(n5833), .Y(n5905) );
  NAND2X0_RVT U5290 ( .A1(n5953), .A2(n5894), .Y(n5833) );
  NAND2X0_RVT U5291 ( .A1(n5773), .A2(n5338), .Y(n5951) );
  INVX0_RVT U5292 ( .A(n5894), .Y(n5773) );
  NAND2X0_RVT U5293 ( .A1(n5660), .A2(n5954), .Y(n5894) );
  AND2X1_RVT U5294 ( .A1(n965), .A2(n974), .Y(n5660) );
  NAND3X0_RVT U5295 ( .A1(n5955), .A2(n5956), .A3(n5957), .Y(n4816) );
  NAND2X0_RVT U5296 ( .A1(n5958), .A2(n5397), .Y(n5957) );
  NAND2X0_RVT U5297 ( .A1(n5959), .A2(n4998), .Y(n5956) );
  NAND2X0_RVT U5298 ( .A1(n5960), .A2(n5961), .Y(n5955) );
  NAND3X0_RVT U5299 ( .A1(n5962), .A2(n5963), .A3(n5403), .Y(n5960) );
  NAND2X0_RVT U5300 ( .A1(n5964), .A2(n5404), .Y(n5963) );
  NAND2X0_RVT U5301 ( .A1(n5832), .A2(n5407), .Y(n5962) );
  NAND3X0_RVT U5302 ( .A1(n5965), .A2(n5966), .A3(n5967), .Y(n4815) );
  NAND2X0_RVT U5303 ( .A1(n5958), .A2(n5411), .Y(n5967) );
  NAND2X0_RVT U5304 ( .A1(n5959), .A2(n5005), .Y(n5966) );
  NAND2X0_RVT U5305 ( .A1(n5968), .A2(n5961), .Y(n5965) );
  NAND3X0_RVT U5306 ( .A1(n5969), .A2(n5970), .A3(n5415), .Y(n5968) );
  NAND2X0_RVT U5307 ( .A1(n5964), .A2(n5416), .Y(n5970) );
  NAND2X0_RVT U5308 ( .A1(n5832), .A2(n5417), .Y(n5969) );
  NAND3X0_RVT U5309 ( .A1(n5971), .A2(n5972), .A3(n5973), .Y(n4814) );
  NAND2X0_RVT U5310 ( .A1(n5958), .A2(n5421), .Y(n5973) );
  NAND2X0_RVT U5311 ( .A1(n5959), .A2(n5012), .Y(n5972) );
  NAND2X0_RVT U5312 ( .A1(n5974), .A2(n5961), .Y(n5971) );
  NAND3X0_RVT U5313 ( .A1(n5975), .A2(n5976), .A3(n5425), .Y(n5974) );
  NAND2X0_RVT U5314 ( .A1(n5964), .A2(n5426), .Y(n5976) );
  NAND2X0_RVT U5315 ( .A1(n5832), .A2(n5427), .Y(n5975) );
  NAND3X0_RVT U5316 ( .A1(n5977), .A2(n5978), .A3(n5979), .Y(n4813) );
  NAND2X0_RVT U5317 ( .A1(n5958), .A2(n5431), .Y(n5979) );
  NAND2X0_RVT U5318 ( .A1(n5959), .A2(n5018), .Y(n5978) );
  NAND2X0_RVT U5319 ( .A1(n5980), .A2(n5961), .Y(n5977) );
  NAND3X0_RVT U5320 ( .A1(n5981), .A2(n5982), .A3(n5435), .Y(n5980) );
  NAND2X0_RVT U5321 ( .A1(n5964), .A2(n5436), .Y(n5982) );
  NAND2X0_RVT U5322 ( .A1(n5832), .A2(n5437), .Y(n5981) );
  NAND3X0_RVT U5323 ( .A1(n5983), .A2(n5984), .A3(n5985), .Y(n4812) );
  NAND2X0_RVT U5324 ( .A1(n5958), .A2(n5441), .Y(n5985) );
  NAND2X0_RVT U5325 ( .A1(n5959), .A2(n5025), .Y(n5984) );
  NAND2X0_RVT U5326 ( .A1(n5986), .A2(n5961), .Y(n5983) );
  NAND3X0_RVT U5327 ( .A1(n5987), .A2(n5988), .A3(n5445), .Y(n5986) );
  NAND2X0_RVT U5328 ( .A1(n5964), .A2(n5446), .Y(n5988) );
  NAND2X0_RVT U5329 ( .A1(n5832), .A2(n5447), .Y(n5987) );
  NAND3X0_RVT U5330 ( .A1(n5989), .A2(n5990), .A3(n5991), .Y(n4811) );
  NAND2X0_RVT U5331 ( .A1(n5958), .A2(n5451), .Y(n5991) );
  NAND2X0_RVT U5332 ( .A1(n5959), .A2(n5032), .Y(n5990) );
  NAND2X0_RVT U5333 ( .A1(n5992), .A2(n5961), .Y(n5989) );
  NAND3X0_RVT U5334 ( .A1(n5993), .A2(n5994), .A3(n5455), .Y(n5992) );
  NAND2X0_RVT U5335 ( .A1(n5964), .A2(n5456), .Y(n5994) );
  NAND2X0_RVT U5336 ( .A1(n5832), .A2(n5457), .Y(n5993) );
  NAND3X0_RVT U5337 ( .A1(n5995), .A2(n5996), .A3(n5997), .Y(n4810) );
  NAND2X0_RVT U5338 ( .A1(n5958), .A2(n5461), .Y(n5997) );
  NAND2X0_RVT U5339 ( .A1(n5959), .A2(n5039), .Y(n5996) );
  NAND2X0_RVT U5340 ( .A1(n5998), .A2(n5961), .Y(n5995) );
  NAND3X0_RVT U5341 ( .A1(n5999), .A2(n6000), .A3(n5465), .Y(n5998) );
  NAND2X0_RVT U5342 ( .A1(n5964), .A2(n5466), .Y(n6000) );
  NAND2X0_RVT U5343 ( .A1(n5832), .A2(n5467), .Y(n5999) );
  NAND3X0_RVT U5344 ( .A1(n6001), .A2(n6002), .A3(n6003), .Y(n4809) );
  NAND2X0_RVT U5345 ( .A1(n5958), .A2(n5329), .Y(n6003) );
  AND2X1_RVT U5346 ( .A1(n5890), .A2(n5961), .Y(n5958) );
  NAND2X0_RVT U5347 ( .A1(n5959), .A2(n5044), .Y(n6002) );
  INVX0_RVT U5348 ( .A(n5961), .Y(n5959) );
  NAND2X0_RVT U5349 ( .A1(n6004), .A2(n5961), .Y(n6001) );
  NAND3X0_RVT U5350 ( .A1(n6005), .A2(n6006), .A3(n6007), .Y(n5961) );
  NAND2X0_RVT U5351 ( .A1(n6008), .A2(n5359), .Y(n6007) );
  NAND2X0_RVT U5352 ( .A1(n5476), .A2(n5891), .Y(n6006) );
  NAND2X0_RVT U5353 ( .A1(n6009), .A2(n5479), .Y(n6005) );
  NAND3X0_RVT U5354 ( .A1(n6010), .A2(n6011), .A3(n5334), .Y(n6004) );
  NAND2X0_RVT U5355 ( .A1(n5964), .A2(n5335), .Y(n6011) );
  INVX0_RVT U5356 ( .A(n5891), .Y(n5964) );
  NAND2X0_RVT U5357 ( .A1(n6012), .A2(n5953), .Y(n5891) );
  NAND2X0_RVT U5358 ( .A1(n5832), .A2(n5338), .Y(n6010) );
  INVX0_RVT U5359 ( .A(n5953), .Y(n5832) );
  NAND2X0_RVT U5360 ( .A1(n5778), .A2(n5895), .Y(n5953) );
  NAND3X0_RVT U5361 ( .A1(n6013), .A2(n6014), .A3(n6015), .Y(n4808) );
  NAND2X0_RVT U5362 ( .A1(n6016), .A2(n5397), .Y(n6015) );
  NAND2X0_RVT U5363 ( .A1(n6017), .A2(n4999), .Y(n6014) );
  NAND2X0_RVT U5364 ( .A1(n6018), .A2(n6019), .Y(n6013) );
  NAND3X0_RVT U5365 ( .A1(n6020), .A2(n6021), .A3(n5403), .Y(n6018) );
  NAND2X0_RVT U5366 ( .A1(n6022), .A2(n5404), .Y(n6021) );
  NAND2X0_RVT U5367 ( .A1(n5890), .A2(n5407), .Y(n6020) );
  NAND3X0_RVT U5368 ( .A1(n6023), .A2(n6024), .A3(n6025), .Y(n4807) );
  NAND2X0_RVT U5369 ( .A1(n6016), .A2(n5411), .Y(n6025) );
  NAND2X0_RVT U5370 ( .A1(n6017), .A2(n5006), .Y(n6024) );
  NAND2X0_RVT U5371 ( .A1(n6026), .A2(n6019), .Y(n6023) );
  NAND3X0_RVT U5372 ( .A1(n6027), .A2(n6028), .A3(n5415), .Y(n6026) );
  NAND2X0_RVT U5373 ( .A1(n6022), .A2(n5416), .Y(n6028) );
  NAND2X0_RVT U5374 ( .A1(n5890), .A2(n5417), .Y(n6027) );
  NAND3X0_RVT U5375 ( .A1(n6029), .A2(n6030), .A3(n6031), .Y(n4806) );
  NAND2X0_RVT U5376 ( .A1(n6016), .A2(n5421), .Y(n6031) );
  NAND2X0_RVT U5377 ( .A1(n6017), .A2(n5013), .Y(n6030) );
  NAND2X0_RVT U5378 ( .A1(n6032), .A2(n6019), .Y(n6029) );
  NAND3X0_RVT U5379 ( .A1(n6033), .A2(n6034), .A3(n5425), .Y(n6032) );
  NAND2X0_RVT U5380 ( .A1(n6022), .A2(n5426), .Y(n6034) );
  NAND2X0_RVT U5381 ( .A1(n5890), .A2(n5427), .Y(n6033) );
  NAND3X0_RVT U5382 ( .A1(n6035), .A2(n6036), .A3(n6037), .Y(n4805) );
  NAND2X0_RVT U5383 ( .A1(n6016), .A2(n5431), .Y(n6037) );
  NAND2X0_RVT U5384 ( .A1(n6017), .A2(n5019), .Y(n6036) );
  NAND2X0_RVT U5385 ( .A1(n6038), .A2(n6019), .Y(n6035) );
  NAND3X0_RVT U5386 ( .A1(n6039), .A2(n6040), .A3(n5435), .Y(n6038) );
  NAND2X0_RVT U5387 ( .A1(n6022), .A2(n5436), .Y(n6040) );
  NAND2X0_RVT U5388 ( .A1(n5890), .A2(n5437), .Y(n6039) );
  NAND3X0_RVT U5389 ( .A1(n6041), .A2(n6042), .A3(n6043), .Y(n4804) );
  NAND2X0_RVT U5390 ( .A1(n6016), .A2(n5441), .Y(n6043) );
  NAND2X0_RVT U5391 ( .A1(n6017), .A2(n5026), .Y(n6042) );
  NAND2X0_RVT U5392 ( .A1(n6044), .A2(n6019), .Y(n6041) );
  NAND3X0_RVT U5393 ( .A1(n6045), .A2(n6046), .A3(n5445), .Y(n6044) );
  NAND2X0_RVT U5394 ( .A1(n6022), .A2(n5446), .Y(n6046) );
  NAND2X0_RVT U5395 ( .A1(n5890), .A2(n5447), .Y(n6045) );
  NAND3X0_RVT U5396 ( .A1(n6047), .A2(n6048), .A3(n6049), .Y(n4803) );
  NAND2X0_RVT U5397 ( .A1(n6016), .A2(n5451), .Y(n6049) );
  NAND2X0_RVT U5398 ( .A1(n6017), .A2(n5033), .Y(n6048) );
  NAND2X0_RVT U5399 ( .A1(n6050), .A2(n6019), .Y(n6047) );
  NAND3X0_RVT U5400 ( .A1(n6051), .A2(n6052), .A3(n5455), .Y(n6050) );
  NAND2X0_RVT U5401 ( .A1(n6022), .A2(n5456), .Y(n6052) );
  NAND2X0_RVT U5402 ( .A1(n5890), .A2(n5457), .Y(n6051) );
  NAND3X0_RVT U5403 ( .A1(n6053), .A2(n6054), .A3(n6055), .Y(n4802) );
  NAND2X0_RVT U5404 ( .A1(n6016), .A2(n5461), .Y(n6055) );
  NAND2X0_RVT U5405 ( .A1(n6017), .A2(n5040), .Y(n6054) );
  NAND2X0_RVT U5406 ( .A1(n6056), .A2(n6019), .Y(n6053) );
  NAND3X0_RVT U5407 ( .A1(n6057), .A2(n6058), .A3(n5465), .Y(n6056) );
  NAND2X0_RVT U5408 ( .A1(n6022), .A2(n5466), .Y(n6058) );
  NAND2X0_RVT U5409 ( .A1(n5890), .A2(n5467), .Y(n6057) );
  NAND3X0_RVT U5410 ( .A1(n6059), .A2(n6060), .A3(n6061), .Y(n4801) );
  NAND2X0_RVT U5411 ( .A1(n6016), .A2(n5329), .Y(n6061) );
  AND2X1_RVT U5412 ( .A1(n5949), .A2(n6019), .Y(n6016) );
  NAND2X0_RVT U5413 ( .A1(n6017), .A2(n5047), .Y(n6060) );
  INVX0_RVT U5414 ( .A(n6019), .Y(n6017) );
  NAND2X0_RVT U5415 ( .A1(n6062), .A2(n6019), .Y(n6059) );
  NAND3X0_RVT U5416 ( .A1(n6063), .A2(n6064), .A3(n6065), .Y(n6019) );
  NAND2X0_RVT U5417 ( .A1(n6066), .A2(n5359), .Y(n6065) );
  NAND2X0_RVT U5418 ( .A1(n5476), .A2(n5950), .Y(n6064) );
  NAND2X0_RVT U5419 ( .A1(n6067), .A2(n5479), .Y(n6063) );
  NAND3X0_RVT U5420 ( .A1(n6068), .A2(n6069), .A3(n5334), .Y(n6062) );
  NAND2X0_RVT U5421 ( .A1(n6022), .A2(n5335), .Y(n6069) );
  INVX0_RVT U5422 ( .A(n5950), .Y(n6022) );
  NAND2X0_RVT U5423 ( .A1(n6070), .A2(n6012), .Y(n5950) );
  NAND2X0_RVT U5424 ( .A1(n5890), .A2(n5338), .Y(n6068) );
  INVX0_RVT U5425 ( .A(n6012), .Y(n5890) );
  NAND2X0_RVT U5426 ( .A1(n5778), .A2(n5954), .Y(n6012) );
  AND2X1_RVT U5427 ( .A1(n965), .A2(n4909), .Y(n5778) );
  NAND3X0_RVT U5428 ( .A1(n6071), .A2(n6072), .A3(n6073), .Y(n4800) );
  NAND2X0_RVT U5429 ( .A1(n6074), .A2(n5397), .Y(n6073) );
  NAND2X0_RVT U5430 ( .A1(n6075), .A2(n5001), .Y(n6072) );
  NAND2X0_RVT U5431 ( .A1(n6076), .A2(n6077), .Y(n6071) );
  NAND3X0_RVT U5432 ( .A1(n6078), .A2(n6079), .A3(n5403), .Y(n6076) );
  NAND2X0_RVT U5433 ( .A1(n6080), .A2(n5404), .Y(n6079) );
  NAND2X0_RVT U5434 ( .A1(n5949), .A2(n5407), .Y(n6078) );
  NAND3X0_RVT U5435 ( .A1(n6081), .A2(n6082), .A3(n6083), .Y(n4799) );
  NAND2X0_RVT U5436 ( .A1(n6074), .A2(n5411), .Y(n6083) );
  NAND2X0_RVT U5437 ( .A1(n6075), .A2(n5008), .Y(n6082) );
  NAND2X0_RVT U5438 ( .A1(n6084), .A2(n6077), .Y(n6081) );
  NAND3X0_RVT U5439 ( .A1(n6085), .A2(n6086), .A3(n5415), .Y(n6084) );
  NAND2X0_RVT U5440 ( .A1(n6080), .A2(n5416), .Y(n6086) );
  NAND2X0_RVT U5441 ( .A1(n5949), .A2(n5417), .Y(n6085) );
  NAND3X0_RVT U5442 ( .A1(n6087), .A2(n6088), .A3(n6089), .Y(n4798) );
  NAND2X0_RVT U5443 ( .A1(n6074), .A2(n5421), .Y(n6089) );
  NAND2X0_RVT U5444 ( .A1(n6075), .A2(n5015), .Y(n6088) );
  NAND2X0_RVT U5445 ( .A1(n6090), .A2(n6077), .Y(n6087) );
  NAND3X0_RVT U5446 ( .A1(n6091), .A2(n6092), .A3(n5425), .Y(n6090) );
  NAND2X0_RVT U5447 ( .A1(n6080), .A2(n5426), .Y(n6092) );
  NAND2X0_RVT U5448 ( .A1(n5949), .A2(n5427), .Y(n6091) );
  NAND3X0_RVT U5449 ( .A1(n6093), .A2(n6094), .A3(n6095), .Y(n4797) );
  NAND2X0_RVT U5450 ( .A1(n6074), .A2(n5431), .Y(n6095) );
  NAND2X0_RVT U5451 ( .A1(n6075), .A2(n5021), .Y(n6094) );
  NAND2X0_RVT U5452 ( .A1(n6096), .A2(n6077), .Y(n6093) );
  NAND3X0_RVT U5453 ( .A1(n6097), .A2(n6098), .A3(n5435), .Y(n6096) );
  NAND2X0_RVT U5454 ( .A1(n6080), .A2(n5436), .Y(n6098) );
  NAND2X0_RVT U5455 ( .A1(n5949), .A2(n5437), .Y(n6097) );
  NAND3X0_RVT U5456 ( .A1(n6099), .A2(n6100), .A3(n6101), .Y(n4796) );
  NAND2X0_RVT U5457 ( .A1(n6074), .A2(n5441), .Y(n6101) );
  NAND2X0_RVT U5458 ( .A1(n6075), .A2(n5028), .Y(n6100) );
  NAND2X0_RVT U5459 ( .A1(n6102), .A2(n6077), .Y(n6099) );
  NAND3X0_RVT U5460 ( .A1(n6103), .A2(n6104), .A3(n5445), .Y(n6102) );
  NAND2X0_RVT U5461 ( .A1(n6080), .A2(n5446), .Y(n6104) );
  NAND2X0_RVT U5462 ( .A1(n5949), .A2(n5447), .Y(n6103) );
  NAND3X0_RVT U5463 ( .A1(n6105), .A2(n6106), .A3(n6107), .Y(n4795) );
  NAND2X0_RVT U5464 ( .A1(n6074), .A2(n5451), .Y(n6107) );
  NAND2X0_RVT U5465 ( .A1(n6075), .A2(n5035), .Y(n6106) );
  NAND2X0_RVT U5466 ( .A1(n6108), .A2(n6077), .Y(n6105) );
  NAND3X0_RVT U5467 ( .A1(n6109), .A2(n6110), .A3(n5455), .Y(n6108) );
  NAND2X0_RVT U5468 ( .A1(n6080), .A2(n5456), .Y(n6110) );
  NAND2X0_RVT U5469 ( .A1(n5949), .A2(n5457), .Y(n6109) );
  NAND3X0_RVT U5470 ( .A1(n6111), .A2(n6112), .A3(n6113), .Y(n4794) );
  NAND2X0_RVT U5471 ( .A1(n6074), .A2(n5461), .Y(n6113) );
  NAND2X0_RVT U5472 ( .A1(n6075), .A2(n5042), .Y(n6112) );
  NAND2X0_RVT U5473 ( .A1(n6114), .A2(n6077), .Y(n6111) );
  NAND3X0_RVT U5474 ( .A1(n6115), .A2(n6116), .A3(n5465), .Y(n6114) );
  NAND2X0_RVT U5475 ( .A1(n6080), .A2(n5466), .Y(n6116) );
  NAND2X0_RVT U5476 ( .A1(n5949), .A2(n5467), .Y(n6115) );
  NAND3X0_RVT U5477 ( .A1(n6117), .A2(n6118), .A3(n6119), .Y(n4793) );
  NAND2X0_RVT U5478 ( .A1(n6074), .A2(n5329), .Y(n6119) );
  AND2X1_RVT U5479 ( .A1(n6008), .A2(n6077), .Y(n6074) );
  NAND2X0_RVT U5480 ( .A1(n6075), .A2(n5051), .Y(n6118) );
  INVX0_RVT U5481 ( .A(n6077), .Y(n6075) );
  NAND2X0_RVT U5482 ( .A1(n6120), .A2(n6077), .Y(n6117) );
  NAND3X0_RVT U5483 ( .A1(n6121), .A2(n6122), .A3(n6123), .Y(n6077) );
  NAND2X0_RVT U5484 ( .A1(n6124), .A2(n5359), .Y(n6123) );
  NAND2X0_RVT U5485 ( .A1(n5476), .A2(n6009), .Y(n6122) );
  NAND2X0_RVT U5486 ( .A1(n6125), .A2(n5479), .Y(n6121) );
  NAND3X0_RVT U5487 ( .A1(n6126), .A2(n6127), .A3(n5334), .Y(n6120) );
  NAND2X0_RVT U5488 ( .A1(n6080), .A2(n5335), .Y(n6127) );
  INVX0_RVT U5489 ( .A(n6009), .Y(n6080) );
  NAND2X0_RVT U5490 ( .A1(n6128), .A2(n6070), .Y(n6009) );
  NAND2X0_RVT U5491 ( .A1(n5949), .A2(n5338), .Y(n6126) );
  INVX0_RVT U5492 ( .A(n6070), .Y(n5949) );
  NAND2X0_RVT U5493 ( .A1(n5659), .A2(n6129), .Y(n6070) );
  NAND3X0_RVT U5494 ( .A1(n6130), .A2(n6131), .A3(n6132), .Y(n4792) );
  NAND2X0_RVT U5495 ( .A1(n6133), .A2(n5397), .Y(n6132) );
  NAND2X0_RVT U5496 ( .A1(n6134), .A2(n5133), .Y(n6131) );
  NAND2X0_RVT U5497 ( .A1(n6135), .A2(n6136), .Y(n6130) );
  NAND3X0_RVT U5498 ( .A1(n6137), .A2(n6138), .A3(n5403), .Y(n6135) );
  NAND2X0_RVT U5499 ( .A1(n6139), .A2(n5404), .Y(n6138) );
  NAND2X0_RVT U5500 ( .A1(n6008), .A2(n5407), .Y(n6137) );
  NAND3X0_RVT U5501 ( .A1(n6140), .A2(n6141), .A3(n6142), .Y(n4791) );
  NAND2X0_RVT U5502 ( .A1(n6133), .A2(n5411), .Y(n6142) );
  NAND2X0_RVT U5503 ( .A1(n6134), .A2(n5138), .Y(n6141) );
  NAND2X0_RVT U5504 ( .A1(n6143), .A2(n6136), .Y(n6140) );
  NAND3X0_RVT U5505 ( .A1(n6144), .A2(n6145), .A3(n5415), .Y(n6143) );
  NAND2X0_RVT U5506 ( .A1(n6139), .A2(n5416), .Y(n6145) );
  NAND2X0_RVT U5507 ( .A1(n6008), .A2(n5417), .Y(n6144) );
  NAND3X0_RVT U5508 ( .A1(n6146), .A2(n6147), .A3(n6148), .Y(n4790) );
  NAND2X0_RVT U5509 ( .A1(n6133), .A2(n5421), .Y(n6148) );
  NAND2X0_RVT U5510 ( .A1(n6134), .A2(n5143), .Y(n6147) );
  NAND2X0_RVT U5511 ( .A1(n6149), .A2(n6136), .Y(n6146) );
  NAND3X0_RVT U5512 ( .A1(n6150), .A2(n6151), .A3(n5425), .Y(n6149) );
  NAND2X0_RVT U5513 ( .A1(n6139), .A2(n5426), .Y(n6151) );
  NAND2X0_RVT U5514 ( .A1(n6008), .A2(n5427), .Y(n6150) );
  NAND3X0_RVT U5515 ( .A1(n6152), .A2(n6153), .A3(n6154), .Y(n4789) );
  NAND2X0_RVT U5516 ( .A1(n6133), .A2(n5431), .Y(n6154) );
  NAND2X0_RVT U5517 ( .A1(n6134), .A2(n5148), .Y(n6153) );
  NAND2X0_RVT U5518 ( .A1(n6155), .A2(n6136), .Y(n6152) );
  NAND3X0_RVT U5519 ( .A1(n6156), .A2(n6157), .A3(n5435), .Y(n6155) );
  NAND2X0_RVT U5520 ( .A1(n6139), .A2(n5436), .Y(n6157) );
  NAND2X0_RVT U5521 ( .A1(n6008), .A2(n5437), .Y(n6156) );
  NAND3X0_RVT U5522 ( .A1(n6158), .A2(n6159), .A3(n6160), .Y(n4788) );
  NAND2X0_RVT U5523 ( .A1(n6133), .A2(n5441), .Y(n6160) );
  NAND2X0_RVT U5524 ( .A1(n6134), .A2(n5153), .Y(n6159) );
  NAND2X0_RVT U5525 ( .A1(n6161), .A2(n6136), .Y(n6158) );
  NAND3X0_RVT U5526 ( .A1(n6162), .A2(n6163), .A3(n5445), .Y(n6161) );
  NAND2X0_RVT U5527 ( .A1(n6139), .A2(n5446), .Y(n6163) );
  NAND2X0_RVT U5528 ( .A1(n6008), .A2(n5447), .Y(n6162) );
  NAND3X0_RVT U5529 ( .A1(n6164), .A2(n6165), .A3(n6166), .Y(n4787) );
  NAND2X0_RVT U5530 ( .A1(n6133), .A2(n5451), .Y(n6166) );
  NAND2X0_RVT U5531 ( .A1(n6134), .A2(n5158), .Y(n6165) );
  NAND2X0_RVT U5532 ( .A1(n6167), .A2(n6136), .Y(n6164) );
  NAND3X0_RVT U5533 ( .A1(n6168), .A2(n6169), .A3(n5455), .Y(n6167) );
  NAND2X0_RVT U5534 ( .A1(n6139), .A2(n5456), .Y(n6169) );
  NAND2X0_RVT U5535 ( .A1(n6008), .A2(n5457), .Y(n6168) );
  NAND3X0_RVT U5536 ( .A1(n6170), .A2(n6171), .A3(n6172), .Y(n4786) );
  NAND2X0_RVT U5537 ( .A1(n6133), .A2(n5461), .Y(n6172) );
  NAND2X0_RVT U5538 ( .A1(n6134), .A2(n5163), .Y(n6171) );
  NAND2X0_RVT U5539 ( .A1(n6173), .A2(n6136), .Y(n6170) );
  NAND3X0_RVT U5540 ( .A1(n6174), .A2(n6175), .A3(n5465), .Y(n6173) );
  NAND2X0_RVT U5541 ( .A1(n6139), .A2(n5466), .Y(n6175) );
  NAND2X0_RVT U5542 ( .A1(n6008), .A2(n5467), .Y(n6174) );
  NAND3X0_RVT U5543 ( .A1(n6176), .A2(n6177), .A3(n6178), .Y(n4785) );
  NAND2X0_RVT U5544 ( .A1(n6133), .A2(n5329), .Y(n6178) );
  AND2X1_RVT U5545 ( .A1(n6066), .A2(n6136), .Y(n6133) );
  NAND2X0_RVT U5546 ( .A1(n6134), .A2(n5171), .Y(n6177) );
  INVX0_RVT U5547 ( .A(n6136), .Y(n6134) );
  NAND2X0_RVT U5548 ( .A1(n6179), .A2(n6136), .Y(n6176) );
  NAND3X0_RVT U5549 ( .A1(n6180), .A2(n6181), .A3(n6182), .Y(n6136) );
  NAND2X0_RVT U5550 ( .A1(n5337), .A2(n5359), .Y(n6182) );
  NAND2X0_RVT U5551 ( .A1(n5476), .A2(n6067), .Y(n6181) );
  NAND2X0_RVT U5552 ( .A1(n6183), .A2(n5479), .Y(n6180) );
  NAND3X0_RVT U5553 ( .A1(n6184), .A2(n6185), .A3(n5334), .Y(n6179) );
  NAND2X0_RVT U5554 ( .A1(n6139), .A2(n5335), .Y(n6185) );
  INVX0_RVT U5555 ( .A(n6067), .Y(n6139) );
  NAND2X0_RVT U5556 ( .A1(n6186), .A2(n6128), .Y(n6067) );
  NAND2X0_RVT U5557 ( .A1(n6008), .A2(n5338), .Y(n6184) );
  INVX0_RVT U5558 ( .A(n6128), .Y(n6008) );
  NAND2X0_RVT U5559 ( .A1(n5719), .A2(n6129), .Y(n6128) );
  NAND3X0_RVT U5560 ( .A1(n6187), .A2(n6188), .A3(n6189), .Y(n4784) );
  NAND2X0_RVT U5561 ( .A1(n6190), .A2(n5397), .Y(n6189) );
  NAND2X0_RVT U5562 ( .A1(n6191), .A2(n4996), .Y(n6188) );
  NAND2X0_RVT U5563 ( .A1(n6192), .A2(n6193), .Y(n6187) );
  NAND3X0_RVT U5564 ( .A1(n6194), .A2(n6195), .A3(n5403), .Y(n6192) );
  NAND2X0_RVT U5565 ( .A1(n6196), .A2(n5404), .Y(n6195) );
  NAND2X0_RVT U5566 ( .A1(n6066), .A2(n5407), .Y(n6194) );
  NAND3X0_RVT U5567 ( .A1(n6197), .A2(n6198), .A3(n6199), .Y(n4783) );
  NAND2X0_RVT U5568 ( .A1(n6190), .A2(n5411), .Y(n6199) );
  NAND2X0_RVT U5569 ( .A1(n6191), .A2(n5003), .Y(n6198) );
  NAND2X0_RVT U5570 ( .A1(n6200), .A2(n6193), .Y(n6197) );
  NAND3X0_RVT U5571 ( .A1(n6201), .A2(n6202), .A3(n5415), .Y(n6200) );
  NAND2X0_RVT U5572 ( .A1(n6196), .A2(n5416), .Y(n6202) );
  NAND2X0_RVT U5573 ( .A1(n6066), .A2(n5417), .Y(n6201) );
  NAND3X0_RVT U5574 ( .A1(n6203), .A2(n6204), .A3(n6205), .Y(n4782) );
  NAND2X0_RVT U5575 ( .A1(n6190), .A2(n5421), .Y(n6205) );
  NAND2X0_RVT U5576 ( .A1(n6191), .A2(n5010), .Y(n6204) );
  NAND2X0_RVT U5577 ( .A1(n6206), .A2(n6193), .Y(n6203) );
  NAND3X0_RVT U5578 ( .A1(n6207), .A2(n6208), .A3(n5425), .Y(n6206) );
  NAND2X0_RVT U5579 ( .A1(n6196), .A2(n5426), .Y(n6208) );
  NAND2X0_RVT U5580 ( .A1(n6066), .A2(n5427), .Y(n6207) );
  NAND3X0_RVT U5581 ( .A1(n6209), .A2(n6210), .A3(n6211), .Y(n4781) );
  NAND2X0_RVT U5582 ( .A1(n6190), .A2(n5431), .Y(n6211) );
  NAND2X0_RVT U5583 ( .A1(n6191), .A2(n5016), .Y(n6210) );
  NAND2X0_RVT U5584 ( .A1(n6212), .A2(n6193), .Y(n6209) );
  NAND3X0_RVT U5585 ( .A1(n6213), .A2(n6214), .A3(n5435), .Y(n6212) );
  NAND2X0_RVT U5586 ( .A1(n6196), .A2(n5436), .Y(n6214) );
  NAND2X0_RVT U5587 ( .A1(n6066), .A2(n5437), .Y(n6213) );
  NAND3X0_RVT U5588 ( .A1(n6215), .A2(n6216), .A3(n6217), .Y(n4780) );
  NAND2X0_RVT U5589 ( .A1(n6190), .A2(n5441), .Y(n6217) );
  NAND2X0_RVT U5590 ( .A1(n6191), .A2(n5023), .Y(n6216) );
  NAND2X0_RVT U5591 ( .A1(n6218), .A2(n6193), .Y(n6215) );
  NAND3X0_RVT U5592 ( .A1(n6219), .A2(n6220), .A3(n5445), .Y(n6218) );
  NAND2X0_RVT U5593 ( .A1(n6196), .A2(n5446), .Y(n6220) );
  NAND2X0_RVT U5594 ( .A1(n6066), .A2(n5447), .Y(n6219) );
  NAND3X0_RVT U5595 ( .A1(n6221), .A2(n6222), .A3(n6223), .Y(n4779) );
  NAND2X0_RVT U5596 ( .A1(n6190), .A2(n5451), .Y(n6223) );
  NAND2X0_RVT U5597 ( .A1(n6191), .A2(n5030), .Y(n6222) );
  NAND2X0_RVT U5598 ( .A1(n6224), .A2(n6193), .Y(n6221) );
  NAND3X0_RVT U5599 ( .A1(n6225), .A2(n6226), .A3(n5455), .Y(n6224) );
  NAND2X0_RVT U5600 ( .A1(n6196), .A2(n5456), .Y(n6226) );
  NAND2X0_RVT U5601 ( .A1(n6066), .A2(n5457), .Y(n6225) );
  NAND3X0_RVT U5602 ( .A1(n6227), .A2(n6228), .A3(n6229), .Y(n4778) );
  NAND2X0_RVT U5603 ( .A1(n6190), .A2(n5461), .Y(n6229) );
  NAND2X0_RVT U5604 ( .A1(n6191), .A2(n5037), .Y(n6228) );
  NAND2X0_RVT U5605 ( .A1(n6230), .A2(n6193), .Y(n6227) );
  NAND3X0_RVT U5606 ( .A1(n6231), .A2(n6232), .A3(n5465), .Y(n6230) );
  NAND2X0_RVT U5607 ( .A1(n6196), .A2(n5466), .Y(n6232) );
  NAND2X0_RVT U5608 ( .A1(n6066), .A2(n5467), .Y(n6231) );
  NAND3X0_RVT U5609 ( .A1(n6233), .A2(n6234), .A3(n6235), .Y(n4777) );
  NAND2X0_RVT U5610 ( .A1(n6190), .A2(n5329), .Y(n6235) );
  AND2X1_RVT U5611 ( .A1(n6124), .A2(n6193), .Y(n6190) );
  NAND2X0_RVT U5612 ( .A1(n6191), .A2(n5045), .Y(n6234) );
  INVX0_RVT U5613 ( .A(n6193), .Y(n6191) );
  NAND2X0_RVT U5614 ( .A1(n6236), .A2(n6193), .Y(n6233) );
  NAND3X0_RVT U5615 ( .A1(n6237), .A2(n6238), .A3(n6239), .Y(n6193) );
  NAND2X0_RVT U5616 ( .A1(n5406), .A2(n5359), .Y(n6239) );
  NAND2X0_RVT U5617 ( .A1(n5476), .A2(n6125), .Y(n6238) );
  NAND2X0_RVT U5618 ( .A1(n6240), .A2(n5479), .Y(n6237) );
  NAND3X0_RVT U5619 ( .A1(n6241), .A2(n6242), .A3(n5334), .Y(n6236) );
  NAND2X0_RVT U5620 ( .A1(n6196), .A2(n5335), .Y(n6242) );
  INVX0_RVT U5621 ( .A(n6125), .Y(n6196) );
  NAND2X0_RVT U5622 ( .A1(n6243), .A2(n6186), .Y(n6125) );
  NAND2X0_RVT U5623 ( .A1(n6066), .A2(n5338), .Y(n6241) );
  INVX0_RVT U5624 ( .A(n6186), .Y(n6066) );
  NAND2X0_RVT U5625 ( .A1(n5659), .A2(n6244), .Y(n6186) );
  AND2X1_RVT U5626 ( .A1(n973), .A2(n975), .Y(n5659) );
  NAND3X0_RVT U5627 ( .A1(n6245), .A2(n6246), .A3(n6247), .Y(n4776) );
  NAND2X0_RVT U5628 ( .A1(n6248), .A2(n5397), .Y(n6247) );
  NAND2X0_RVT U5629 ( .A1(n6249), .A2(n5117), .Y(n6246) );
  NAND2X0_RVT U5630 ( .A1(n6250), .A2(n6251), .Y(n6245) );
  NAND3X0_RVT U5631 ( .A1(n6252), .A2(n6253), .A3(n5403), .Y(n6250) );
  NAND2X0_RVT U5632 ( .A1(n6254), .A2(n5404), .Y(n6253) );
  NAND2X0_RVT U5633 ( .A1(n6124), .A2(n5407), .Y(n6252) );
  NAND3X0_RVT U5634 ( .A1(n6255), .A2(n6256), .A3(n6257), .Y(n4775) );
  NAND2X0_RVT U5635 ( .A1(n6248), .A2(n5411), .Y(n6257) );
  NAND2X0_RVT U5636 ( .A1(n6249), .A2(n5112), .Y(n6256) );
  NAND2X0_RVT U5637 ( .A1(n6258), .A2(n6251), .Y(n6255) );
  NAND3X0_RVT U5638 ( .A1(n6259), .A2(n6260), .A3(n5415), .Y(n6258) );
  NAND2X0_RVT U5639 ( .A1(n6254), .A2(n5416), .Y(n6260) );
  NAND2X0_RVT U5640 ( .A1(n6124), .A2(n5417), .Y(n6259) );
  NAND3X0_RVT U5641 ( .A1(n6261), .A2(n6262), .A3(n6263), .Y(n4774) );
  NAND2X0_RVT U5642 ( .A1(n6248), .A2(n5421), .Y(n6263) );
  NAND2X0_RVT U5643 ( .A1(n6249), .A2(n5113), .Y(n6262) );
  NAND2X0_RVT U5644 ( .A1(n6264), .A2(n6251), .Y(n6261) );
  NAND3X0_RVT U5645 ( .A1(n6265), .A2(n6266), .A3(n5425), .Y(n6264) );
  NAND2X0_RVT U5646 ( .A1(n6254), .A2(n5426), .Y(n6266) );
  NAND2X0_RVT U5647 ( .A1(n6124), .A2(n5427), .Y(n6265) );
  NAND3X0_RVT U5648 ( .A1(n6267), .A2(n6268), .A3(n6269), .Y(n4773) );
  NAND2X0_RVT U5649 ( .A1(n6248), .A2(n5431), .Y(n6269) );
  NAND2X0_RVT U5650 ( .A1(n6249), .A2(n5114), .Y(n6268) );
  NAND2X0_RVT U5651 ( .A1(n6270), .A2(n6251), .Y(n6267) );
  NAND3X0_RVT U5652 ( .A1(n6271), .A2(n6272), .A3(n5435), .Y(n6270) );
  NAND2X0_RVT U5653 ( .A1(n6254), .A2(n5436), .Y(n6272) );
  NAND2X0_RVT U5654 ( .A1(n6124), .A2(n5437), .Y(n6271) );
  NAND3X0_RVT U5655 ( .A1(n6273), .A2(n6274), .A3(n6275), .Y(n4772) );
  NAND2X0_RVT U5656 ( .A1(n6248), .A2(n5441), .Y(n6275) );
  NAND2X0_RVT U5657 ( .A1(n6249), .A2(n5115), .Y(n6274) );
  NAND2X0_RVT U5658 ( .A1(n6276), .A2(n6251), .Y(n6273) );
  NAND3X0_RVT U5659 ( .A1(n6277), .A2(n6278), .A3(n5445), .Y(n6276) );
  NAND2X0_RVT U5660 ( .A1(n6254), .A2(n5446), .Y(n6278) );
  NAND2X0_RVT U5661 ( .A1(n6124), .A2(n5447), .Y(n6277) );
  NAND3X0_RVT U5662 ( .A1(n6279), .A2(n6280), .A3(n6281), .Y(n4771) );
  NAND2X0_RVT U5663 ( .A1(n6248), .A2(n5451), .Y(n6281) );
  NAND2X0_RVT U5664 ( .A1(n6249), .A2(n5116), .Y(n6280) );
  NAND2X0_RVT U5665 ( .A1(n6282), .A2(n6251), .Y(n6279) );
  NAND3X0_RVT U5666 ( .A1(n6283), .A2(n6284), .A3(n5455), .Y(n6282) );
  NAND2X0_RVT U5667 ( .A1(n6254), .A2(n5456), .Y(n6284) );
  NAND2X0_RVT U5668 ( .A1(n6124), .A2(n5457), .Y(n6283) );
  NAND3X0_RVT U5669 ( .A1(n6285), .A2(n6286), .A3(n6287), .Y(n4770) );
  NAND2X0_RVT U5670 ( .A1(n6248), .A2(n5461), .Y(n6287) );
  NAND2X0_RVT U5671 ( .A1(n6249), .A2(n5111), .Y(n6286) );
  NAND2X0_RVT U5672 ( .A1(n6288), .A2(n6251), .Y(n6285) );
  NAND3X0_RVT U5673 ( .A1(n6289), .A2(n6290), .A3(n5465), .Y(n6288) );
  NAND2X0_RVT U5674 ( .A1(n6254), .A2(n5466), .Y(n6290) );
  NAND2X0_RVT U5675 ( .A1(n6124), .A2(n5467), .Y(n6289) );
  NAND3X0_RVT U5676 ( .A1(n6291), .A2(n6292), .A3(n6293), .Y(n4769) );
  NAND2X0_RVT U5677 ( .A1(n6248), .A2(n5329), .Y(n6293) );
  XNOR2X1_RVT U5678 ( .A1(n6294), .A2(Datai[23]), .Y(n5329) );
  NAND2X0_RVT U5679 ( .A1(Datai[22]), .A2(n6295), .Y(n6294) );
  AND2X1_RVT U5680 ( .A1(n5337), .A2(n6251), .Y(n6248) );
  NAND2X0_RVT U5681 ( .A1(n6249), .A2(n5048), .Y(n6292) );
  INVX0_RVT U5682 ( .A(n6251), .Y(n6249) );
  NAND2X0_RVT U5683 ( .A1(n6296), .A2(n6251), .Y(n6291) );
  NAND3X0_RVT U5684 ( .A1(n6297), .A2(n6298), .A3(n6299), .Y(n6251) );
  NAND2X0_RVT U5685 ( .A1(n5471), .A2(n5359), .Y(n6299) );
  INVX0_RVT U5686 ( .A(n6300), .Y(n5471) );
  NAND2X0_RVT U5687 ( .A1(n5476), .A2(n6183), .Y(n6298) );
  NAND2X0_RVT U5688 ( .A1(n5477), .A2(n5479), .Y(n6297) );
  NAND2X0_RVT U5689 ( .A1(n6301), .A2(n6300), .Y(n5477) );
  NAND3X0_RVT U5690 ( .A1(n6302), .A2(n6303), .A3(n5334), .Y(n6296) );
  AND2X1_RVT U5691 ( .A1(n6304), .A2(n6305), .Y(n5334) );
  NAND2X0_RVT U5692 ( .A1(n6306), .A2(n6307), .Y(n6305) );
  NAND2X0_RVT U5693 ( .A1(Datai[7]), .A2(n6308), .Y(n6304) );
  NAND2X0_RVT U5694 ( .A1(n6254), .A2(n5335), .Y(n6303) );
  AND2X1_RVT U5695 ( .A1(Datai[7]), .A2(n5371), .Y(n5335) );
  INVX0_RVT U5696 ( .A(n6183), .Y(n6254) );
  NAND2X0_RVT U5697 ( .A1(n6309), .A2(n6243), .Y(n6183) );
  NAND2X0_RVT U5698 ( .A1(n6124), .A2(n5338), .Y(n6302) );
  AND2X1_RVT U5699 ( .A1(n6310), .A2(n6311), .Y(n5338) );
  NAND2X0_RVT U5700 ( .A1(Datai[30]), .A2(n6312), .Y(n6311) );
  INVX0_RVT U5701 ( .A(n6243), .Y(n6124) );
  NAND2X0_RVT U5702 ( .A1(n5719), .A2(n6244), .Y(n6243) );
  AND2X1_RVT U5703 ( .A1(n973), .A2(n4928), .Y(n5719) );
  NAND3X0_RVT U5704 ( .A1(n6313), .A2(n6314), .A3(n6315), .Y(n4768) );
  NAND2X0_RVT U5705 ( .A1(n5328), .A2(n5397), .Y(n6315) );
  OR2X1_RVT U5706 ( .A1(n5330), .A2(n815), .Y(n6314) );
  NAND2X0_RVT U5707 ( .A1(n6316), .A2(n5330), .Y(n6313) );
  NAND3X0_RVT U5708 ( .A1(n6317), .A2(n6318), .A3(n5403), .Y(n6316) );
  AND2X1_RVT U5709 ( .A1(n6319), .A2(n6320), .Y(n5403) );
  NAND2X0_RVT U5710 ( .A1(n6306), .A2(n6321), .Y(n6320) );
  NAND2X0_RVT U5711 ( .A1(Datai[0]), .A2(n6308), .Y(n6319) );
  NAND2X0_RVT U5712 ( .A1(n5404), .A2(n5336), .Y(n6318) );
  AND2X1_RVT U5713 ( .A1(Datai[0]), .A2(n5371), .Y(n5404) );
  NAND2X0_RVT U5714 ( .A1(n5337), .A2(n5407), .Y(n6317) );
  NAND3X0_RVT U5715 ( .A1(n6322), .A2(n6323), .A3(n6324), .Y(n4767) );
  NAND2X0_RVT U5716 ( .A1(n5328), .A2(n5411), .Y(n6324) );
  OR2X1_RVT U5717 ( .A1(n5330), .A2(n813), .Y(n6323) );
  NAND2X0_RVT U5718 ( .A1(n6325), .A2(n5330), .Y(n6322) );
  NAND3X0_RVT U5719 ( .A1(n6326), .A2(n6327), .A3(n5415), .Y(n6325) );
  AND2X1_RVT U5720 ( .A1(n6328), .A2(n6329), .Y(n5415) );
  NAND2X0_RVT U5721 ( .A1(n6306), .A2(n6330), .Y(n6329) );
  NAND2X0_RVT U5722 ( .A1(Datai[1]), .A2(n6308), .Y(n6328) );
  NAND2X0_RVT U5723 ( .A1(n5416), .A2(n5336), .Y(n6327) );
  AND2X1_RVT U5724 ( .A1(Datai[1]), .A2(n5371), .Y(n5416) );
  NAND2X0_RVT U5725 ( .A1(n5337), .A2(n5417), .Y(n6326) );
  NAND3X0_RVT U5726 ( .A1(n6331), .A2(n6332), .A3(n6333), .Y(n4766) );
  NAND2X0_RVT U5727 ( .A1(n5421), .A2(n5328), .Y(n6333) );
  OR2X1_RVT U5728 ( .A1(n5330), .A2(n811), .Y(n6332) );
  NAND2X0_RVT U5729 ( .A1(n6334), .A2(n5330), .Y(n6331) );
  NAND3X0_RVT U5730 ( .A1(n6335), .A2(n6336), .A3(n5425), .Y(n6334) );
  AND2X1_RVT U5731 ( .A1(n6337), .A2(n6338), .Y(n5425) );
  NAND2X0_RVT U5732 ( .A1(n6306), .A2(n6339), .Y(n6338) );
  NAND2X0_RVT U5733 ( .A1(Datai[2]), .A2(n6308), .Y(n6337) );
  NAND2X0_RVT U5734 ( .A1(n5426), .A2(n5336), .Y(n6336) );
  AND2X1_RVT U5735 ( .A1(Datai[2]), .A2(n5371), .Y(n5426) );
  NAND2X0_RVT U5736 ( .A1(n5337), .A2(n5427), .Y(n6335) );
  NAND3X0_RVT U5737 ( .A1(n6340), .A2(n6341), .A3(n6342), .Y(n4765) );
  NAND2X0_RVT U5738 ( .A1(n5431), .A2(n5328), .Y(n6342) );
  OR2X1_RVT U5739 ( .A1(n5330), .A2(n809), .Y(n6341) );
  NAND2X0_RVT U5740 ( .A1(n6343), .A2(n5330), .Y(n6340) );
  NAND3X0_RVT U5741 ( .A1(n6344), .A2(n6345), .A3(n5435), .Y(n6343) );
  AND2X1_RVT U5742 ( .A1(n6346), .A2(n6347), .Y(n5435) );
  NAND2X0_RVT U5743 ( .A1(n6306), .A2(n6348), .Y(n6347) );
  NAND2X0_RVT U5744 ( .A1(Datai[3]), .A2(n6308), .Y(n6346) );
  NAND2X0_RVT U5745 ( .A1(n5436), .A2(n5336), .Y(n6345) );
  AND2X1_RVT U5746 ( .A1(Datai[3]), .A2(n5371), .Y(n5436) );
  NAND2X0_RVT U5747 ( .A1(n5337), .A2(n5437), .Y(n6344) );
  NAND3X0_RVT U5748 ( .A1(n6349), .A2(n6350), .A3(n6351), .Y(n4764) );
  NAND2X0_RVT U5749 ( .A1(n5441), .A2(n5328), .Y(n6351) );
  XNOR2X1_RVT U5750 ( .A1(n6352), .A2(Datai[20]), .Y(n5441) );
  OR2X1_RVT U5751 ( .A1(n5330), .A2(n807), .Y(n6350) );
  NAND2X0_RVT U5752 ( .A1(n6353), .A2(n5330), .Y(n6349) );
  NAND3X0_RVT U5753 ( .A1(n6354), .A2(n6355), .A3(n5445), .Y(n6353) );
  AND2X1_RVT U5754 ( .A1(n6356), .A2(n6357), .Y(n5445) );
  NAND2X0_RVT U5755 ( .A1(n6306), .A2(n6358), .Y(n6357) );
  NAND2X0_RVT U5756 ( .A1(Datai[4]), .A2(n6308), .Y(n6356) );
  NAND2X0_RVT U5757 ( .A1(n5446), .A2(n5336), .Y(n6355) );
  AND2X1_RVT U5758 ( .A1(Datai[4]), .A2(n5371), .Y(n5446) );
  NAND2X0_RVT U5759 ( .A1(n5447), .A2(n5337), .Y(n6354) );
  XOR2X1_RVT U5760 ( .A1(n6359), .A2(n6360), .Y(n5447) );
  NAND3X0_RVT U5761 ( .A1(n6361), .A2(n6362), .A3(n6363), .Y(n4763) );
  NAND2X0_RVT U5762 ( .A1(n5451), .A2(n5328), .Y(n6363) );
  XOR2X1_RVT U5763 ( .A1(n6364), .A2(Datai[21]), .Y(n5451) );
  OR2X1_RVT U5764 ( .A1(n5330), .A2(n805), .Y(n6362) );
  NAND2X0_RVT U5765 ( .A1(n6365), .A2(n5330), .Y(n6361) );
  NAND3X0_RVT U5766 ( .A1(n6366), .A2(n6367), .A3(n5455), .Y(n6365) );
  AND2X1_RVT U5767 ( .A1(n6368), .A2(n6369), .Y(n5455) );
  NAND2X0_RVT U5768 ( .A1(n6306), .A2(n6370), .Y(n6369) );
  NAND2X0_RVT U5769 ( .A1(Datai[5]), .A2(n6308), .Y(n6368) );
  NAND2X0_RVT U5770 ( .A1(n5456), .A2(n5336), .Y(n6367) );
  AND2X1_RVT U5771 ( .A1(Datai[5]), .A2(n5371), .Y(n5456) );
  NAND2X0_RVT U5772 ( .A1(n5337), .A2(n5457), .Y(n6366) );
  XOR2X1_RVT U5773 ( .A1(Datai[29]), .A2(n6371), .Y(n5457) );
  NAND3X0_RVT U5774 ( .A1(n6372), .A2(n6373), .A3(n6374), .Y(n4762) );
  NAND2X0_RVT U5775 ( .A1(n5328), .A2(n5461), .Y(n6374) );
  XOR2X1_RVT U5776 ( .A1(n6295), .A2(Datai[22]), .Y(n5461) );
  AND2X1_RVT U5777 ( .A1(Datai[21]), .A2(n6364), .Y(n6295) );
  NOR2X0_RVT U5778 ( .A1(n6375), .A2(n6352), .Y(n6364) );
  NAND2X0_RVT U5779 ( .A1(n6376), .A2(n6377), .Y(n6352) );
  INVX0_RVT U5780 ( .A(n6378), .Y(n6376) );
  AND2X1_RVT U5781 ( .A1(n5406), .A2(n5330), .Y(n5328) );
  INVX0_RVT U5782 ( .A(n6301), .Y(n5406) );
  OR2X1_RVT U5783 ( .A1(n5330), .A2(n803), .Y(n6373) );
  NAND2X0_RVT U5784 ( .A1(n6379), .A2(n5330), .Y(n6372) );
  NAND2X0_RVT U5785 ( .A1(n5359), .A2(n5532), .Y(n6382) );
  INVX0_RVT U5786 ( .A(n5599), .Y(n5532) );
  NAND2X0_RVT U5787 ( .A1(n5476), .A2(n6240), .Y(n6381) );
  NAND2X0_RVT U5788 ( .A1(n5537), .A2(n5479), .Y(n6380) );
  NAND2X0_RVT U5789 ( .A1(n5599), .A2(n6300), .Y(n5537) );
  NAND2X0_RVT U5790 ( .A1(n6244), .A2(n5895), .Y(n6300) );
  NAND2X0_RVT U5791 ( .A1(n6244), .A2(n5954), .Y(n5599) );
  AND2X1_RVT U5792 ( .A1(n4909), .A2(n4930), .Y(n6244) );
  NAND3X0_RVT U5793 ( .A1(n6383), .A2(n6384), .A3(n5465), .Y(n6379) );
  AND2X1_RVT U5794 ( .A1(n6385), .A2(n6386), .Y(n5465) );
  NAND2X0_RVT U5795 ( .A1(n6306), .A2(n6387), .Y(n6386) );
  NAND2X0_RVT U5796 ( .A1(Datai[6]), .A2(n6308), .Y(n6385) );
  NAND2X0_RVT U5797 ( .A1(n5466), .A2(n5336), .Y(n6384) );
  INVX0_RVT U5798 ( .A(n6240), .Y(n5336) );
  NAND2X0_RVT U5799 ( .A1(n6301), .A2(n6309), .Y(n6240) );
  NAND2X0_RVT U5800 ( .A1(n5954), .A2(n6129), .Y(n6301) );
  AND2X1_RVT U5801 ( .A1(n4928), .A2(n4907), .Y(n5954) );
  AND2X1_RVT U5802 ( .A1(Datai[6]), .A2(n5371), .Y(n5466) );
  NAND2X0_RVT U5803 ( .A1(n5337), .A2(n5467), .Y(n6383) );
  INVX0_RVT U5804 ( .A(n6309), .Y(n5337) );
  NAND2X0_RVT U5805 ( .A1(n5895), .A2(n6129), .Y(n6309) );
  AND2X1_RVT U5806 ( .A1(n974), .A2(n4930), .Y(n6129) );
  AND2X1_RVT U5807 ( .A1(n975), .A2(n4907), .Y(n5895) );
  NAND2X0_RVT U5808 ( .A1(n6388), .A2(n6389), .Y(n4761) );
  NAND2X0_RVT U5809 ( .A1(n6390), .A2(n4908), .Y(n6389) );
  NAND2X0_RVT U5810 ( .A1(n6391), .A2(n6392), .Y(n6390) );
  NAND2X0_RVT U5811 ( .A1(n6393), .A2(n5265), .Y(n6392) );
  NAND2X0_RVT U5812 ( .A1(n6394), .A2(n6391), .Y(n6388) );
  NAND3X0_RVT U5813 ( .A1(n6395), .A2(n6396), .A3(n6397), .Y(n6394) );
  NAND2X0_RVT U5814 ( .A1(n5357), .A2(n976), .Y(n6397) );
  NAND3X0_RVT U5815 ( .A1(n939), .A2(n6398), .A3(n5265), .Y(n6396) );
  NAND2X0_RVT U5816 ( .A1(n5359), .A2(n5397), .Y(n6395) );
  NAND2X0_RVT U5817 ( .A1(n6399), .A2(n6400), .Y(n4760) );
  NAND2X0_RVT U5818 ( .A1(n6401), .A2(n6391), .Y(n6400) );
  NAND2X0_RVT U5819 ( .A1(n6402), .A2(n6403), .Y(n6401) );
  NAND3X0_RVT U5820 ( .A1(n936), .A2(n6404), .A3(n5265), .Y(n6403) );
  INVX0_RVT U5821 ( .A(n5431), .Y(n6402) );
  NAND2X0_RVT U5822 ( .A1(n6405), .A2(n4906), .Y(n6399) );
  NAND2X0_RVT U5823 ( .A1(n6391), .A2(n6406), .Y(n6405) );
  OR2X1_RVT U5824 ( .A1(n6404), .A2(n6407), .Y(n6406) );
  NAND2X0_RVT U5825 ( .A1(n6408), .A2(n6409), .Y(n4759) );
  NAND2X0_RVT U5826 ( .A1(n5324), .A2(n4926), .Y(n6409) );
  NAND2X0_RVT U5827 ( .A1(n6410), .A2(n6391), .Y(n6408) );
  NAND3X0_RVT U5828 ( .A1(n6411), .A2(n6412), .A3(n6413), .Y(n6410) );
  NAND2X0_RVT U5829 ( .A1(n5421), .A2(n5359), .Y(n6413) );
  NAND3X0_RVT U5830 ( .A1(n6414), .A2(n4931), .A3(n5357), .Y(n6412) );
  NAND2X0_RVT U5831 ( .A1(n6415), .A2(n6416), .Y(n4758) );
  NAND2X0_RVT U5832 ( .A1(n5324), .A2(n4927), .Y(n6416) );
  INVX0_RVT U5833 ( .A(n6391), .Y(n5324) );
  NAND2X0_RVT U5834 ( .A1(n6417), .A2(n6391), .Y(n6415) );
  NAND3X0_RVT U5835 ( .A1(n5382), .A2(n5340), .A3(n6418), .Y(n6391) );
  NAND3X0_RVT U5836 ( .A1(n6419), .A2(n6420), .A3(n6421), .Y(n6417) );
  NAND2X0_RVT U5837 ( .A1(n5359), .A2(n5411), .Y(n6421) );
  OR3X1_RVT U5838 ( .A1(n5339), .A2(n976), .A3(n6414), .Y(n6420) );
  XNOR2X1_RVT U5839 ( .A1(n9575), .A2(n6422), .Y(n6414) );
  NAND2X0_RVT U5840 ( .A1(n5265), .A2(n6423), .Y(n6419) );
  NAND2X0_RVT U5841 ( .A1(n6424), .A2(n6425), .Y(n4757) );
  NAND2X0_RVT U5842 ( .A1(n5342), .A2(n4969), .Y(n6425) );
  NAND2X0_RVT U5843 ( .A1(n6426), .A2(n6427), .Y(n6424) );
  NAND4X0_RVT U5844 ( .A1(n5380), .A2(n6428), .A3(n6429), .A4(n6430), .Y(n6426) );
  AND4X1_RVT U5845 ( .A1(n6431), .A2(n6432), .A3(n6433), .A4(n6434), .Y(n6430)
         );
  NAND2X0_RVT U5846 ( .A1(READY_n), .A2(n6435), .Y(n6431) );
  NAND2X0_RVT U5847 ( .A1(n6436), .A2(n5263), .Y(n6435) );
  NAND2X0_RVT U5848 ( .A1(n5358), .A2(n5357), .Y(n6428) );
  NAND4X0_RVT U5849 ( .A1(n6437), .A2(n5390), .A3(n6438), .A4(n6439), .Y(n4756) );
  AND3X1_RVT U5850 ( .A1(n6432), .A2(n6407), .A3(n5368), .Y(n6439) );
  NAND2X0_RVT U5851 ( .A1(n6440), .A2(n5268), .Y(n6438) );
  NAND2X0_RVT U5852 ( .A1(n5342), .A2(n4905), .Y(n6437) );
  NAND2X0_RVT U5853 ( .A1(n6441), .A2(n6442), .Y(n4755) );
  NAND2X0_RVT U5854 ( .A1(n5342), .A2(n4910), .Y(n6442) );
  INVX0_RVT U5855 ( .A(n6427), .Y(n5342) );
  NAND2X0_RVT U5856 ( .A1(n6443), .A2(n6427), .Y(n6441) );
  NAND4X0_RVT U5857 ( .A1(n5261), .A2(n5264), .A3(n6429), .A4(n6444), .Y(n6427) );
  AND3X1_RVT U5858 ( .A1(n5340), .A2(n6445), .A3(n5339), .Y(n6444) );
  AND2X1_RVT U5859 ( .A1(n6446), .A2(n6447), .Y(n6429) );
  NAND2X0_RVT U5860 ( .A1(n5265), .A2(n6448), .Y(n6447) );
  NAND4X0_RVT U5861 ( .A1(n5358), .A2(n6449), .A3(n6450), .A4(n6451), .Y(n6448) );
  AND3X1_RVT U5862 ( .A1(n6452), .A2(n6453), .A3(n6454), .Y(n6451) );
  NAND2X0_RVT U5863 ( .A1(n6455), .A2(n6456), .Y(n6454) );
  NAND2X0_RVT U5864 ( .A1(n9513), .A2(n9561), .Y(n6456) );
  INVX0_RVT U5865 ( .A(n6457), .Y(n6455) );
  NAND2X0_RVT U5866 ( .A1(n6458), .A2(n6459), .Y(n6452) );
  NAND2X0_RVT U5867 ( .A1(n6460), .A2(n6461), .Y(n6459) );
  NAND2X0_RVT U5868 ( .A1(n6462), .A2(n6463), .Y(n6461) );
  NAND3X0_RVT U5869 ( .A1(n6464), .A2(n6465), .A3(n6466), .Y(n6463) );
  NAND2X0_RVT U5870 ( .A1(n973), .A2(n6467), .Y(n6466) );
  NAND2X0_RVT U5871 ( .A1(n974), .A2(n6468), .Y(n6465) );
  OR2X1_RVT U5872 ( .A1(n6469), .A2(n6423), .Y(n6468) );
  NAND2X0_RVT U5873 ( .A1(n6423), .A2(n6469), .Y(n6464) );
  NAND2X0_RVT U5874 ( .A1(n6470), .A2(n4928), .Y(n6469) );
  XNOR2X1_RVT U5875 ( .A1(n939), .A2(n6393), .Y(n6470) );
  INVX0_RVT U5876 ( .A(n6398), .Y(n6393) );
  XNOR3X1_RVT U5877 ( .A1(n938), .A2(n6471), .A3(n6472), .Y(n6423) );
  OR2X1_RVT U5878 ( .A1(n6467), .A2(n973), .Y(n6462) );
  NAND2X0_RVT U5879 ( .A1(n965), .A2(n6473), .Y(n6460) );
  OR2X1_RVT U5880 ( .A1(n6473), .A2(n965), .Y(n6458) );
  INVX0_RVT U5881 ( .A(n6474), .Y(n6450) );
  NAND2X0_RVT U5882 ( .A1(n6475), .A2(n6476), .Y(n6449) );
  INVX0_RVT U5883 ( .A(n5383), .Y(n5358) );
  NAND2X0_RVT U5884 ( .A1(n6477), .A2(n6478), .Y(n5383) );
  NAND2X0_RVT U5885 ( .A1(n6479), .A2(n6480), .Y(n6478) );
  NAND2X0_RVT U5886 ( .A1(n6481), .A2(n6482), .Y(n6480) );
  NAND2X0_RVT U5887 ( .A1(n6483), .A2(n5265), .Y(n6482) );
  NAND2X0_RVT U5888 ( .A1(n6483), .A2(n6484), .Y(n6481) );
  NAND2X0_RVT U5889 ( .A1(n5407), .A2(n5417), .Y(n6484) );
  NAND2X0_RVT U5890 ( .A1(n6485), .A2(n6486), .Y(n5417) );
  NAND2X0_RVT U5891 ( .A1(n938), .A2(n6487), .Y(n6486) );
  XNOR2X1_RVT U5892 ( .A1(n6488), .A2(n6489), .Y(n6485) );
  XNOR2X1_RVT U5893 ( .A1(n6490), .A2(n6491), .Y(n5407) );
  NAND2X0_RVT U5894 ( .A1(Datai[24]), .A2(n6492), .Y(n6490) );
  INVX0_RVT U5895 ( .A(n5427), .Y(n6483) );
  NAND2X0_RVT U5896 ( .A1(n6493), .A2(n6494), .Y(n5427) );
  NAND3X0_RVT U5897 ( .A1(n6411), .A2(n6487), .A3(n6495), .Y(n6494) );
  NAND2X0_RVT U5898 ( .A1(n6496), .A2(n4926), .Y(n6495) );
  NAND2X0_RVT U5899 ( .A1(n5265), .A2(n6467), .Y(n6411) );
  XNOR3X1_RVT U5900 ( .A1(n937), .A2(n6497), .A3(n6498), .Y(n6467) );
  XNOR2X1_RVT U5901 ( .A1(n6499), .A2(n6500), .Y(n6493) );
  INVX0_RVT U5902 ( .A(n5437), .Y(n6479) );
  NAND2X0_RVT U5903 ( .A1(n6501), .A2(n6502), .Y(n5437) );
  NAND3X0_RVT U5904 ( .A1(n6503), .A2(n6487), .A3(n936), .Y(n6502) );
  NAND2X0_RVT U5905 ( .A1(n6473), .A2(n5265), .Y(n6503) );
  XNOR2X1_RVT U5906 ( .A1(n6404), .A2(n936), .Y(n6473) );
  NAND2X0_RVT U5907 ( .A1(n6504), .A2(n6505), .Y(n6404) );
  NAND2X0_RVT U5908 ( .A1(n6506), .A2(n4926), .Y(n6505) );
  NAND2X0_RVT U5909 ( .A1(n6498), .A2(n6497), .Y(n6506) );
  OR2X1_RVT U5910 ( .A1(n6498), .A2(n6497), .Y(n6504) );
  NAND2X0_RVT U5911 ( .A1(n6507), .A2(n4927), .Y(n6498) );
  NAND2X0_RVT U5912 ( .A1(n6472), .A2(n6471), .Y(n6507) );
  NAND2X0_RVT U5913 ( .A1(n4908), .A2(n6398), .Y(n6471) );
  NAND2X0_RVT U5914 ( .A1(n6497), .A2(n6508), .Y(n6398) );
  NAND2X0_RVT U5915 ( .A1(n6509), .A2(n6510), .Y(n6508) );
  XNOR2X1_RVT U5916 ( .A1(n6511), .A2(n6512), .Y(n6501) );
  INVX0_RVT U5917 ( .A(n5467), .Y(n6477) );
  XOR2X1_RVT U5918 ( .A1(n6513), .A2(n6312), .Y(n5467) );
  NAND2X0_RVT U5919 ( .A1(n6514), .A2(n6515), .Y(n6312) );
  NAND2X0_RVT U5920 ( .A1(Datai[29]), .A2(n6371), .Y(n6515) );
  NAND2X0_RVT U5921 ( .A1(n6371), .A2(n6487), .Y(n6514) );
  NAND2X0_RVT U5922 ( .A1(n6516), .A2(n6517), .Y(n6371) );
  NAND2X0_RVT U5923 ( .A1(n6360), .A2(n6359), .Y(n6517) );
  AND2X1_RVT U5924 ( .A1(n6511), .A2(n6512), .Y(n6359) );
  OR2X1_RVT U5925 ( .A1(n6487), .A2(Datai[27]), .Y(n6512) );
  AND2X1_RVT U5926 ( .A1(n6499), .A2(n6500), .Y(n6511) );
  OR2X1_RVT U5927 ( .A1(n6487), .A2(Datai[26]), .Y(n6500) );
  AND2X1_RVT U5928 ( .A1(n6488), .A2(n6489), .Y(n6499) );
  NAND2X0_RVT U5929 ( .A1(n6492), .A2(n6518), .Y(n6489) );
  NAND2X0_RVT U5930 ( .A1(Datai[24]), .A2(n6491), .Y(n6518) );
  XNOR2X1_RVT U5931 ( .A1(n6519), .A2(n6492), .Y(n6491) );
  NAND2X0_RVT U5932 ( .A1(n6520), .A2(n6521), .Y(n6519) );
  NAND2X0_RVT U5933 ( .A1(n5476), .A2(n6522), .Y(n6521) );
  NAND2X0_RVT U5934 ( .A1(n6523), .A2(n6524), .Y(n6522) );
  NAND2X0_RVT U5935 ( .A1(Datai[31]), .A2(n6525), .Y(n6524) );
  NAND4X0_RVT U5936 ( .A1(n6526), .A2(n6375), .A3(n6527), .A4(n6528), .Y(n6525) );
  NOR4X0_RVT U5937 ( .A1(n6529), .A2(Datai[16]), .A3(Datai[17]), .A4(Datai[18]), .Y(n6528) );
  NOR3X0_RVT U5938 ( .A1(Datai[22]), .A2(Datai[23]), .A3(Datai[21]), .Y(n6527)
         );
  INVX0_RVT U5939 ( .A(Datai[20]), .Y(n6375) );
  INVX0_RVT U5940 ( .A(Datai[19]), .Y(n6526) );
  NAND2X0_RVT U5941 ( .A1(n6496), .A2(n4908), .Y(n6520) );
  INVX0_RVT U5942 ( .A(n6487), .Y(n6492) );
  OR2X1_RVT U5943 ( .A1(n6487), .A2(Datai[25]), .Y(n6488) );
  AND2X1_RVT U5944 ( .A1(Datai[28]), .A2(n5476), .Y(n6360) );
  AND2X1_RVT U5945 ( .A1(n9561), .A2(n5357), .Y(n6496) );
  OR2X1_RVT U5946 ( .A1(n6487), .A2(Datai[30]), .Y(n6513) );
  NAND2X0_RVT U5947 ( .A1(n6407), .A2(n5339), .Y(n6487) );
  AND3X1_RVT U5948 ( .A1(n6530), .A2(n5263), .A3(n5380), .Y(n5261) );
  NAND2X0_RVT U5949 ( .A1(n5214), .A2(n5268), .Y(n6530) );
  NAND4X0_RVT U5950 ( .A1(n6531), .A2(n6407), .A3(n6532), .A4(n6533), .Y(n6443) );
  OR2X1_RVT U5951 ( .A1(n6436), .A2(READY_n), .Y(n6533) );
  NAND2X0_RVT U5952 ( .A1(n6440), .A2(READY_n), .Y(n6532) );
  INVX0_RVT U5953 ( .A(n5263), .Y(n6440) );
  NAND3X0_RVT U5954 ( .A1(n6534), .A2(n4910), .A3(n790), .Y(n5263) );
  NAND2X0_RVT U5955 ( .A1(n6535), .A2(n6536), .Y(n4754) );
  NAND2X0_RVT U5956 ( .A1(n6537), .A2(n6474), .Y(n6536) );
  NAND2X0_RVT U5957 ( .A1(n6538), .A2(n5110), .Y(n6535) );
  NAND4X0_RVT U5958 ( .A1(n6539), .A2(n6540), .A3(n6541), .A4(n6542), .Y(n4753) );
  NAND2X0_RVT U5959 ( .A1(n5319), .A2(n6543), .Y(n6542) );
  NAND2X0_RVT U5960 ( .A1(n5321), .A2(n6544), .Y(n6541) );
  NAND2X0_RVT U5961 ( .A1(n6545), .A2(n4931), .Y(n6540) );
  NAND4X0_RVT U5962 ( .A1(n6546), .A2(n6547), .A3(n6548), .A4(n6549), .Y(n4752) );
  NAND2X0_RVT U5963 ( .A1(n6550), .A2(n5319), .Y(n6549) );
  NAND2X0_RVT U5964 ( .A1(n5321), .A2(n6551), .Y(n6548) );
  OR2X1_RVT U5965 ( .A1(n5323), .A2(n9568), .Y(n6547) );
  NAND4X0_RVT U5966 ( .A1(n6552), .A2(n6553), .A3(n6554), .A4(n6555), .Y(n4751) );
  NAND2X0_RVT U5967 ( .A1(n6556), .A2(n5319), .Y(n6555) );
  NAND2X0_RVT U5968 ( .A1(n5321), .A2(n6557), .Y(n6554) );
  NAND2X0_RVT U5969 ( .A1(n6545), .A2(n4915), .Y(n6553) );
  NAND4X0_RVT U5970 ( .A1(n6558), .A2(n6559), .A3(n6560), .A4(n6561), .Y(n4750) );
  NAND2X0_RVT U5971 ( .A1(n6562), .A2(n5319), .Y(n6561) );
  NAND2X0_RVT U5972 ( .A1(n5321), .A2(n6563), .Y(n6560) );
  NAND2X0_RVT U5973 ( .A1(n6545), .A2(n4970), .Y(n6559) );
  NAND4X0_RVT U5974 ( .A1(n6564), .A2(n6565), .A3(n6566), .A4(n6567), .Y(n4749) );
  NAND2X0_RVT U5975 ( .A1(n6568), .A2(n5319), .Y(n6567) );
  NAND2X0_RVT U5976 ( .A1(n5321), .A2(n6569), .Y(n6566) );
  NAND2X0_RVT U5977 ( .A1(n6545), .A2(n4916), .Y(n6565) );
  NAND4X0_RVT U5978 ( .A1(n6570), .A2(n6571), .A3(n6572), .A4(n6573), .Y(n4748) );
  NAND2X0_RVT U5979 ( .A1(n6574), .A2(n5319), .Y(n6573) );
  NAND2X0_RVT U5980 ( .A1(n5321), .A2(n6575), .Y(n6572) );
  NAND2X0_RVT U5981 ( .A1(n6545), .A2(n4979), .Y(n6571) );
  NAND4X0_RVT U5982 ( .A1(n6576), .A2(n6577), .A3(n6578), .A4(n6579), .Y(n4747) );
  NAND2X0_RVT U5983 ( .A1(n6580), .A2(n5319), .Y(n6579) );
  NAND2X0_RVT U5984 ( .A1(n5321), .A2(n6581), .Y(n6578) );
  NAND2X0_RVT U5985 ( .A1(n6545), .A2(n4917), .Y(n6577) );
  NAND4X0_RVT U5986 ( .A1(n6582), .A2(n6583), .A3(n6584), .A4(n6585), .Y(n4746) );
  NAND2X0_RVT U5987 ( .A1(n6586), .A2(n5319), .Y(n6585) );
  NAND2X0_RVT U5988 ( .A1(n5321), .A2(n6587), .Y(n6584) );
  NAND2X0_RVT U5989 ( .A1(n6545), .A2(n4971), .Y(n6583) );
  NAND4X0_RVT U5990 ( .A1(n6588), .A2(n6589), .A3(n6590), .A4(n6591), .Y(n4745) );
  NAND2X0_RVT U5991 ( .A1(n6592), .A2(n5319), .Y(n6591) );
  NAND2X0_RVT U5992 ( .A1(n5321), .A2(n6593), .Y(n6590) );
  NAND2X0_RVT U5993 ( .A1(n6545), .A2(n4918), .Y(n6589) );
  NAND4X0_RVT U5994 ( .A1(n6594), .A2(n6595), .A3(n6596), .A4(n6597), .Y(n4744) );
  NAND2X0_RVT U5995 ( .A1(n6598), .A2(n5319), .Y(n6597) );
  NAND2X0_RVT U5996 ( .A1(n5321), .A2(n6599), .Y(n6596) );
  NAND2X0_RVT U5997 ( .A1(n6545), .A2(n4972), .Y(n6595) );
  NAND4X0_RVT U5998 ( .A1(n6600), .A2(n6601), .A3(n6602), .A4(n6603), .Y(n4743) );
  NAND2X0_RVT U5999 ( .A1(n6604), .A2(n5319), .Y(n6603) );
  NAND2X0_RVT U6000 ( .A1(n5321), .A2(n6605), .Y(n6602) );
  NAND2X0_RVT U6001 ( .A1(n6545), .A2(n4919), .Y(n6601) );
  NAND4X0_RVT U6002 ( .A1(n6606), .A2(n6607), .A3(n6608), .A4(n6609), .Y(n4742) );
  NAND2X0_RVT U6003 ( .A1(n6610), .A2(n5319), .Y(n6609) );
  NAND2X0_RVT U6004 ( .A1(n5321), .A2(n6611), .Y(n6608) );
  NAND2X0_RVT U6005 ( .A1(n6545), .A2(n4973), .Y(n6607) );
  NAND4X0_RVT U6006 ( .A1(n6612), .A2(n6613), .A3(n6614), .A4(n6615), .Y(n4741) );
  NAND2X0_RVT U6007 ( .A1(n6616), .A2(n5319), .Y(n6615) );
  NAND2X0_RVT U6008 ( .A1(n5321), .A2(n6617), .Y(n6614) );
  NAND2X0_RVT U6009 ( .A1(n6545), .A2(n4920), .Y(n6613) );
  NAND4X0_RVT U6010 ( .A1(n6618), .A2(n6619), .A3(n6620), .A4(n6621), .Y(n4740) );
  NAND2X0_RVT U6011 ( .A1(n6622), .A2(n5319), .Y(n6621) );
  NAND2X0_RVT U6012 ( .A1(n5321), .A2(n6623), .Y(n6620) );
  NAND2X0_RVT U6013 ( .A1(n6545), .A2(n4974), .Y(n6619) );
  NAND4X0_RVT U6014 ( .A1(n6624), .A2(n6625), .A3(n6626), .A4(n6627), .Y(n4739) );
  NAND2X0_RVT U6015 ( .A1(n6628), .A2(n5319), .Y(n6627) );
  NAND2X0_RVT U6016 ( .A1(n5321), .A2(n6629), .Y(n6626) );
  NAND2X0_RVT U6017 ( .A1(n6545), .A2(n4921), .Y(n6625) );
  NAND4X0_RVT U6018 ( .A1(n6630), .A2(n6631), .A3(n6632), .A4(n6633), .Y(n4738) );
  NAND2X0_RVT U6019 ( .A1(n6634), .A2(n5319), .Y(n6633) );
  NAND2X0_RVT U6020 ( .A1(n5321), .A2(n6635), .Y(n6632) );
  NAND2X0_RVT U6021 ( .A1(n6545), .A2(n4975), .Y(n6631) );
  NAND4X0_RVT U6022 ( .A1(n6636), .A2(n6637), .A3(n6638), .A4(n6639), .Y(n4737) );
  NAND2X0_RVT U6023 ( .A1(n6640), .A2(n5319), .Y(n6639) );
  NAND2X0_RVT U6024 ( .A1(n5321), .A2(n6641), .Y(n6638) );
  NAND2X0_RVT U6025 ( .A1(n6545), .A2(n4922), .Y(n6637) );
  NAND4X0_RVT U6026 ( .A1(n6642), .A2(n6643), .A3(n6644), .A4(n6645), .Y(n4736) );
  NAND2X0_RVT U6027 ( .A1(n6646), .A2(n5319), .Y(n6645) );
  NAND2X0_RVT U6028 ( .A1(n5321), .A2(n6647), .Y(n6644) );
  NAND2X0_RVT U6029 ( .A1(n6545), .A2(n4976), .Y(n6643) );
  NAND4X0_RVT U6030 ( .A1(n6648), .A2(n6649), .A3(n6650), .A4(n6651), .Y(n4735) );
  NAND2X0_RVT U6031 ( .A1(n6652), .A2(n5319), .Y(n6651) );
  NAND2X0_RVT U6032 ( .A1(n5321), .A2(n6653), .Y(n6650) );
  NAND2X0_RVT U6033 ( .A1(n6545), .A2(n4923), .Y(n6649) );
  NAND4X0_RVT U6034 ( .A1(n6654), .A2(n6655), .A3(n6656), .A4(n6657), .Y(n4734) );
  NAND2X0_RVT U6035 ( .A1(n6658), .A2(n5319), .Y(n6657) );
  NAND2X0_RVT U6036 ( .A1(n5321), .A2(n6659), .Y(n6656) );
  NAND2X0_RVT U6037 ( .A1(n6545), .A2(n4977), .Y(n6655) );
  NAND4X0_RVT U6038 ( .A1(n6660), .A2(n6661), .A3(n6662), .A4(n6663), .Y(n4733) );
  NAND2X0_RVT U6039 ( .A1(n6664), .A2(n5319), .Y(n6663) );
  NAND2X0_RVT U6040 ( .A1(n5321), .A2(n6665), .Y(n6662) );
  NAND2X0_RVT U6041 ( .A1(n6545), .A2(n4924), .Y(n6661) );
  NAND4X0_RVT U6042 ( .A1(n6666), .A2(n6667), .A3(n6668), .A4(n6669), .Y(n4732) );
  NAND2X0_RVT U6043 ( .A1(n6670), .A2(n5319), .Y(n6669) );
  NAND2X0_RVT U6044 ( .A1(n5321), .A2(n6671), .Y(n6668) );
  NAND2X0_RVT U6045 ( .A1(n6545), .A2(n4978), .Y(n6667) );
  NAND4X0_RVT U6046 ( .A1(n6672), .A2(n6673), .A3(n6674), .A4(n6675), .Y(n4731) );
  NAND2X0_RVT U6047 ( .A1(n6676), .A2(n5319), .Y(n6675) );
  NAND2X0_RVT U6048 ( .A1(n5321), .A2(n6677), .Y(n6674) );
  NAND2X0_RVT U6049 ( .A1(n6545), .A2(n4965), .Y(n6673) );
  NAND4X0_RVT U6050 ( .A1(n6678), .A2(n6679), .A3(n6680), .A4(n6681), .Y(n4730) );
  NAND2X0_RVT U6051 ( .A1(n5319), .A2(n6682), .Y(n6681) );
  NAND2X0_RVT U6052 ( .A1(n6683), .A2(n5321), .Y(n6680) );
  NAND2X0_RVT U6053 ( .A1(n6545), .A2(n4912), .Y(n6679) );
  NAND4X0_RVT U6054 ( .A1(n6684), .A2(n6685), .A3(n6686), .A4(n6687), .Y(n4729) );
  NAND2X0_RVT U6055 ( .A1(n5319), .A2(n6688), .Y(n6687) );
  NAND2X0_RVT U6056 ( .A1(n6689), .A2(n5321), .Y(n6686) );
  NAND2X0_RVT U6057 ( .A1(n6545), .A2(n5102), .Y(n6685) );
  NAND4X0_RVT U6058 ( .A1(n6690), .A2(n6691), .A3(n6692), .A4(n6693), .Y(n4728) );
  NAND2X0_RVT U6059 ( .A1(n5319), .A2(n6694), .Y(n6693) );
  NAND2X0_RVT U6060 ( .A1(n6695), .A2(n5321), .Y(n6692) );
  NAND2X0_RVT U6061 ( .A1(n6545), .A2(n5103), .Y(n6691) );
  NAND4X0_RVT U6062 ( .A1(n6696), .A2(n6697), .A3(n6698), .A4(n6699), .Y(n4727) );
  NAND2X0_RVT U6063 ( .A1(n5319), .A2(n6700), .Y(n6699) );
  NAND2X0_RVT U6064 ( .A1(n6701), .A2(n5321), .Y(n6698) );
  NAND2X0_RVT U6065 ( .A1(n6545), .A2(n5104), .Y(n6697) );
  NAND4X0_RVT U6066 ( .A1(n6702), .A2(n6703), .A3(n6704), .A4(n6705), .Y(n4726) );
  NAND2X0_RVT U6067 ( .A1(n5319), .A2(n6706), .Y(n6705) );
  NAND2X0_RVT U6068 ( .A1(n6707), .A2(n5321), .Y(n6704) );
  NAND2X0_RVT U6069 ( .A1(n6545), .A2(n5105), .Y(n6703) );
  NAND4X0_RVT U6070 ( .A1(n6708), .A2(n6709), .A3(n6710), .A4(n6711), .Y(n4725) );
  NAND2X0_RVT U6071 ( .A1(n5319), .A2(n6712), .Y(n6711) );
  NAND2X0_RVT U6072 ( .A1(n6713), .A2(n5321), .Y(n6710) );
  NAND2X0_RVT U6073 ( .A1(n6545), .A2(n5106), .Y(n6709) );
  NAND4X0_RVT U6074 ( .A1(n6714), .A2(n6715), .A3(n6716), .A4(n6717), .Y(n4724) );
  NAND2X0_RVT U6075 ( .A1(n6718), .A2(n5319), .Y(n6717) );
  NAND2X0_RVT U6076 ( .A1(n5321), .A2(n6719), .Y(n6716) );
  NAND2X0_RVT U6077 ( .A1(n6545), .A2(n5107), .Y(n6715) );
  NAND4X0_RVT U6078 ( .A1(n6720), .A2(n6721), .A3(n6722), .A4(n6723), .Y(n4723) );
  NAND2X0_RVT U6079 ( .A1(n6724), .A2(n5319), .Y(n6723) );
  NAND3X0_RVT U6080 ( .A1(n6727), .A2(n6728), .A3(n6509), .Y(n6726) );
  NAND2X0_RVT U6081 ( .A1(n5321), .A2(n6729), .Y(n6722) );
  NAND2X0_RVT U6082 ( .A1(n6545), .A2(n5052), .Y(n6721) );
  NAND2X0_RVT U6083 ( .A1(n6731), .A2(n6418), .Y(n5323) );
  NAND2X0_RVT U6084 ( .A1(n5265), .A2(n6732), .Y(n6418) );
  NAND3X0_RVT U6085 ( .A1(n6728), .A2(n6497), .A3(n6472), .Y(n6732) );
  NAND3X0_RVT U6086 ( .A1(n6733), .A2(n6734), .A3(n6735), .Y(n4722) );
  NAND2X0_RVT U6087 ( .A1(n6736), .A2(n6434), .Y(n6735) );
  OR2X1_RVT U6088 ( .A1(n6537), .A2(n9513), .Y(n6734) );
  NAND3X0_RVT U6089 ( .A1(n6475), .A2(n6476), .A3(n6537), .Y(n6733) );
  INVX0_RVT U6090 ( .A(n6538), .Y(n6537) );
  NAND2X0_RVT U6091 ( .A1(n5265), .A2(n6457), .Y(n6538) );
  NAND4X0_RVT U6092 ( .A1(n6737), .A2(n6738), .A3(n6739), .A4(n6740), .Y(n6457) );
  NAND2X0_RVT U6093 ( .A1(n6741), .A2(n5268), .Y(n6740) );
  OR2X1_RVT U6094 ( .A1(n6742), .A2(n5271), .Y(n6741) );
  INVX0_RVT U6095 ( .A(n6730), .Y(n6737) );
  NAND2X0_RVT U6096 ( .A1(n6743), .A2(n6453), .Y(n6730) );
  NAND2X0_RVT U6097 ( .A1(n6744), .A2(n6745), .Y(n4721) );
  OR2X1_RVT U6098 ( .A1(n6746), .A2(n9512), .Y(n6745) );
  NAND2X0_RVT U6099 ( .A1(n6747), .A2(n6746), .Y(n6744) );
  NAND2X0_RVT U6100 ( .A1(n6748), .A2(n5264), .Y(n6747) );
  NAND2X0_RVT U6101 ( .A1(n6749), .A2(n6750), .Y(n4720) );
  NAND2X0_RVT U6102 ( .A1(n5276), .A2(W_R_n), .Y(n6750) );
  NAND2X0_RVT U6103 ( .A1(n9512), .A2(n6751), .Y(n6749) );
  NAND2X0_RVT U6104 ( .A1(n6752), .A2(n6753), .Y(n4719) );
  NAND2X0_RVT U6105 ( .A1(n5260), .A2(n5173), .Y(n6753) );
  INVX0_RVT U6106 ( .A(n6746), .Y(n5260) );
  NAND2X0_RVT U6107 ( .A1(n6754), .A2(n6746), .Y(n6752) );
  NAND2X0_RVT U6108 ( .A1(n5264), .A2(n6755), .Y(n6746) );
  NAND2X0_RVT U6109 ( .A1(n5264), .A2(n6756), .Y(n6754) );
  AND2X1_RVT U6110 ( .A1(n6433), .A2(n6436), .Y(n5264) );
  NAND2X0_RVT U6111 ( .A1(n6757), .A2(n6758), .Y(n4718) );
  NAND2X0_RVT U6112 ( .A1(n5276), .A2(M_IO_n), .Y(n6758) );
  NAND2X0_RVT U6113 ( .A1(n6751), .A2(n5173), .Y(n6757) );
  NAND2X0_RVT U6114 ( .A1(n6436), .A2(n6759), .Y(n4717) );
  NAND2X0_RVT U6115 ( .A1(n6755), .A2(n5195), .Y(n6759) );
  NAND2X0_RVT U6116 ( .A1(n6760), .A2(n6534), .Y(n6436) );
  NAND3X0_RVT U6117 ( .A1(n6761), .A2(n6762), .A3(n5294), .Y(n4716) );
  NAND3X0_RVT U6118 ( .A1(n732), .A2(n731), .A3(n730), .Y(n5294) );
  NAND2X0_RVT U6119 ( .A1(n5276), .A2(D_C_n), .Y(n6762) );
  NAND2X0_RVT U6120 ( .A1(n9511), .A2(n6751), .Y(n6761) );
  NAND4X0_RVT U6121 ( .A1(n6763), .A2(n6764), .A3(n6765), .A4(n6766), .Y(n4715) );
  NAND2X0_RVT U6122 ( .A1(n5203), .A2(n4961), .Y(n6766) );
  NAND2X0_RVT U6123 ( .A1(n6767), .A2(n5211), .Y(n6765) );
  NAND2X0_RVT U6124 ( .A1(n5196), .A2(Datai[0]), .Y(n6764) );
  NAND2X0_RVT U6125 ( .A1(n6769), .A2(n5210), .Y(n6763) );
  NAND4X0_RVT U6126 ( .A1(n6770), .A2(n6771), .A3(n6772), .A4(n6773), .Y(n4714) );
  NAND2X0_RVT U6127 ( .A1(n5202), .A2(n4959), .Y(n6773) );
  NAND2X0_RVT U6128 ( .A1(n6774), .A2(n5209), .Y(n6772) );
  NAND2X0_RVT U6129 ( .A1(n5199), .A2(Datai[1]), .Y(n6771) );
  NAND2X0_RVT U6130 ( .A1(n6775), .A2(n5208), .Y(n6770) );
  NAND4X0_RVT U6131 ( .A1(n6776), .A2(n6777), .A3(n6778), .A4(n6779), .Y(n4713) );
  NAND2X0_RVT U6132 ( .A1(n5201), .A2(n4957), .Y(n6779) );
  NAND2X0_RVT U6133 ( .A1(n6780), .A2(n5211), .Y(n6778) );
  NAND2X0_RVT U6134 ( .A1(n5198), .A2(Datai[2]), .Y(n6777) );
  NAND2X0_RVT U6135 ( .A1(n6781), .A2(n5210), .Y(n6776) );
  NAND4X0_RVT U6136 ( .A1(n6782), .A2(n6783), .A3(n6784), .A4(n6785), .Y(n4712) );
  NAND2X0_RVT U6137 ( .A1(n5200), .A2(n4951), .Y(n6785) );
  NAND2X0_RVT U6138 ( .A1(n6786), .A2(n5209), .Y(n6784) );
  NAND2X0_RVT U6139 ( .A1(n5197), .A2(Datai[3]), .Y(n6783) );
  NAND2X0_RVT U6140 ( .A1(n6787), .A2(n5208), .Y(n6782) );
  NAND4X0_RVT U6141 ( .A1(n6788), .A2(n6789), .A3(n6790), .A4(n6791), .Y(n4711) );
  NAND2X0_RVT U6142 ( .A1(n5203), .A2(n4954), .Y(n6791) );
  NAND2X0_RVT U6143 ( .A1(n6792), .A2(n5211), .Y(n6790) );
  NAND2X0_RVT U6144 ( .A1(n5196), .A2(Datai[4]), .Y(n6789) );
  NAND2X0_RVT U6145 ( .A1(n6793), .A2(n5210), .Y(n6788) );
  NAND4X0_RVT U6146 ( .A1(n6794), .A2(n6795), .A3(n6796), .A4(n6797), .Y(n4710) );
  NAND2X0_RVT U6147 ( .A1(n5202), .A2(n4948), .Y(n6797) );
  NAND2X0_RVT U6148 ( .A1(n6798), .A2(n5209), .Y(n6796) );
  NAND2X0_RVT U6149 ( .A1(n5199), .A2(Datai[5]), .Y(n6795) );
  NAND2X0_RVT U6150 ( .A1(n6799), .A2(n5208), .Y(n6794) );
  NAND4X0_RVT U6151 ( .A1(n6800), .A2(n6801), .A3(n6802), .A4(n6803), .Y(n4709) );
  NAND2X0_RVT U6152 ( .A1(n5201), .A2(n4956), .Y(n6803) );
  NAND2X0_RVT U6153 ( .A1(n6804), .A2(n5211), .Y(n6802) );
  NAND2X0_RVT U6154 ( .A1(n5198), .A2(Datai[6]), .Y(n6801) );
  NAND2X0_RVT U6155 ( .A1(n6805), .A2(n5210), .Y(n6800) );
  NAND4X0_RVT U6156 ( .A1(n6806), .A2(n6807), .A3(n6808), .A4(n6809), .Y(n4708) );
  NAND2X0_RVT U6157 ( .A1(n5200), .A2(n4950), .Y(n6809) );
  NAND2X0_RVT U6158 ( .A1(n6810), .A2(n5209), .Y(n6808) );
  NAND2X0_RVT U6159 ( .A1(n5197), .A2(Datai[7]), .Y(n6807) );
  NAND2X0_RVT U6160 ( .A1(n6811), .A2(n5208), .Y(n6806) );
  NAND4X0_RVT U6161 ( .A1(n6812), .A2(n6813), .A3(n6814), .A4(n6815), .Y(n4707) );
  NAND2X0_RVT U6162 ( .A1(n5203), .A2(n4953), .Y(n6815) );
  NAND2X0_RVT U6163 ( .A1(n6816), .A2(n5211), .Y(n6814) );
  NAND2X0_RVT U6164 ( .A1(Datai[8]), .A2(n5199), .Y(n6813) );
  NAND2X0_RVT U6165 ( .A1(n6817), .A2(n5210), .Y(n6812) );
  NAND4X0_RVT U6166 ( .A1(n6818), .A2(n6819), .A3(n6820), .A4(n6821), .Y(n4706) );
  NAND2X0_RVT U6167 ( .A1(n5202), .A2(n4947), .Y(n6821) );
  NAND2X0_RVT U6168 ( .A1(n6822), .A2(n5209), .Y(n6820) );
  NAND2X0_RVT U6169 ( .A1(Datai[9]), .A2(n5198), .Y(n6819) );
  NAND2X0_RVT U6170 ( .A1(n6823), .A2(n5208), .Y(n6818) );
  NAND4X0_RVT U6171 ( .A1(n6824), .A2(n6825), .A3(n6826), .A4(n6827), .Y(n4705) );
  NAND2X0_RVT U6172 ( .A1(n5201), .A2(n4952), .Y(n6827) );
  NAND2X0_RVT U6173 ( .A1(n6828), .A2(n5211), .Y(n6826) );
  NAND2X0_RVT U6174 ( .A1(Datai[10]), .A2(n5197), .Y(n6825) );
  NAND2X0_RVT U6175 ( .A1(n6829), .A2(n5210), .Y(n6824) );
  NAND4X0_RVT U6176 ( .A1(n6830), .A2(n6831), .A3(n6832), .A4(n6833), .Y(n4704) );
  NAND2X0_RVT U6177 ( .A1(n5200), .A2(n4946), .Y(n6833) );
  NAND2X0_RVT U6178 ( .A1(n6834), .A2(n5209), .Y(n6832) );
  NAND2X0_RVT U6179 ( .A1(Datai[11]), .A2(n5196), .Y(n6831) );
  NAND2X0_RVT U6180 ( .A1(n6835), .A2(n5208), .Y(n6830) );
  NAND4X0_RVT U6181 ( .A1(n6836), .A2(n6837), .A3(n6838), .A4(n6839), .Y(n4703) );
  NAND2X0_RVT U6182 ( .A1(n5203), .A2(n4955), .Y(n6839) );
  NAND2X0_RVT U6183 ( .A1(n6840), .A2(n5211), .Y(n6838) );
  NAND2X0_RVT U6184 ( .A1(Datai[12]), .A2(n5199), .Y(n6837) );
  NAND2X0_RVT U6185 ( .A1(n6841), .A2(n5210), .Y(n6836) );
  NAND4X0_RVT U6186 ( .A1(n6842), .A2(n6843), .A3(n6844), .A4(n6845), .Y(n4702) );
  NAND2X0_RVT U6187 ( .A1(n5202), .A2(n4949), .Y(n6845) );
  NAND2X0_RVT U6188 ( .A1(n6846), .A2(n5209), .Y(n6844) );
  NAND2X0_RVT U6189 ( .A1(Datai[13]), .A2(n5198), .Y(n6843) );
  NAND2X0_RVT U6190 ( .A1(n6847), .A2(n5208), .Y(n6842) );
  NAND4X0_RVT U6191 ( .A1(n6848), .A2(n6849), .A3(n6850), .A4(n6851), .Y(n4701) );
  NAND2X0_RVT U6192 ( .A1(n5201), .A2(n4960), .Y(n6851) );
  NAND2X0_RVT U6193 ( .A1(n6852), .A2(n5211), .Y(n6850) );
  NAND2X0_RVT U6194 ( .A1(Datai[14]), .A2(n5197), .Y(n6849) );
  NAND2X0_RVT U6195 ( .A1(n6853), .A2(n5210), .Y(n6848) );
  NAND4X0_RVT U6196 ( .A1(n6854), .A2(n6855), .A3(n6856), .A4(n6857), .Y(n4700) );
  NAND2X0_RVT U6197 ( .A1(n5200), .A2(n4945), .Y(n6857) );
  NAND2X0_RVT U6198 ( .A1(n6858), .A2(n5209), .Y(n6856) );
  NAND2X0_RVT U6199 ( .A1(Datai[15]), .A2(n5196), .Y(n6855) );
  NAND2X0_RVT U6200 ( .A1(n6859), .A2(n5208), .Y(n6854) );
  NAND3X0_RVT U6201 ( .A1(n6860), .A2(n6861), .A3(n6862), .Y(n4699) );
  NAND2X0_RVT U6202 ( .A1(n6863), .A2(n5176), .Y(n6862) );
  NAND2X0_RVT U6203 ( .A1(n6864), .A2(n4961), .Y(n6860) );
  NAND3X0_RVT U6204 ( .A1(n6865), .A2(n6866), .A3(n6867), .Y(n4698) );
  NAND2X0_RVT U6205 ( .A1(n6863), .A2(n5175), .Y(n6867) );
  NAND2X0_RVT U6206 ( .A1(n6864), .A2(n4959), .Y(n6865) );
  NAND3X0_RVT U6207 ( .A1(n6868), .A2(n6869), .A3(n6870), .Y(n4697) );
  NAND2X0_RVT U6208 ( .A1(n6863), .A2(n5177), .Y(n6870) );
  NAND2X0_RVT U6209 ( .A1(n6864), .A2(n4957), .Y(n6868) );
  NAND3X0_RVT U6210 ( .A1(n6871), .A2(n6872), .A3(n6873), .Y(n4696) );
  NAND2X0_RVT U6211 ( .A1(n6863), .A2(n5178), .Y(n6873) );
  NAND2X0_RVT U6212 ( .A1(n6864), .A2(n4951), .Y(n6871) );
  NAND3X0_RVT U6213 ( .A1(n6874), .A2(n6875), .A3(n6876), .Y(n4695) );
  NAND2X0_RVT U6214 ( .A1(n6863), .A2(n5179), .Y(n6876) );
  NAND2X0_RVT U6215 ( .A1(n6864), .A2(n4954), .Y(n6874) );
  NAND3X0_RVT U6216 ( .A1(n6877), .A2(n6878), .A3(n6879), .Y(n4694) );
  NAND2X0_RVT U6217 ( .A1(n6863), .A2(n5180), .Y(n6879) );
  NAND2X0_RVT U6218 ( .A1(n6864), .A2(n4948), .Y(n6877) );
  NAND3X0_RVT U6219 ( .A1(n6880), .A2(n6881), .A3(n6882), .Y(n4693) );
  NAND2X0_RVT U6220 ( .A1(n6863), .A2(n5181), .Y(n6882) );
  NAND2X0_RVT U6221 ( .A1(n6864), .A2(n4956), .Y(n6880) );
  NAND3X0_RVT U6222 ( .A1(n6883), .A2(n6884), .A3(n6885), .Y(n4692) );
  NAND2X0_RVT U6223 ( .A1(n6863), .A2(n5182), .Y(n6885) );
  NAND2X0_RVT U6224 ( .A1(n6864), .A2(n4950), .Y(n6883) );
  NAND3X0_RVT U6225 ( .A1(n6886), .A2(n6887), .A3(n6888), .Y(n4691) );
  NAND2X0_RVT U6226 ( .A1(n6863), .A2(n5183), .Y(n6888) );
  NAND2X0_RVT U6227 ( .A1(n6864), .A2(n4953), .Y(n6886) );
  NAND3X0_RVT U6228 ( .A1(n6889), .A2(n6890), .A3(n6891), .Y(n4690) );
  NAND2X0_RVT U6229 ( .A1(n6863), .A2(n5184), .Y(n6891) );
  NAND2X0_RVT U6230 ( .A1(n6864), .A2(n4947), .Y(n6889) );
  NAND3X0_RVT U6231 ( .A1(n6892), .A2(n6893), .A3(n6894), .Y(n4689) );
  NAND2X0_RVT U6232 ( .A1(n6863), .A2(n5185), .Y(n6894) );
  NAND2X0_RVT U6233 ( .A1(n6864), .A2(n4952), .Y(n6892) );
  NAND3X0_RVT U6234 ( .A1(n6895), .A2(n6896), .A3(n6897), .Y(n4688) );
  NAND2X0_RVT U6235 ( .A1(n6863), .A2(n5186), .Y(n6897) );
  NAND2X0_RVT U6236 ( .A1(n6864), .A2(n4946), .Y(n6895) );
  NAND3X0_RVT U6237 ( .A1(n6898), .A2(n6899), .A3(n6900), .Y(n4687) );
  NAND2X0_RVT U6238 ( .A1(n6863), .A2(n5187), .Y(n6900) );
  NAND2X0_RVT U6239 ( .A1(n6864), .A2(n4955), .Y(n6898) );
  NAND3X0_RVT U6240 ( .A1(n6901), .A2(n6902), .A3(n6903), .Y(n4686) );
  NAND2X0_RVT U6241 ( .A1(n6863), .A2(n5188), .Y(n6903) );
  NAND2X0_RVT U6242 ( .A1(n6864), .A2(n4949), .Y(n6901) );
  NAND3X0_RVT U6243 ( .A1(n6904), .A2(n6905), .A3(n6906), .Y(n4685) );
  NAND2X0_RVT U6244 ( .A1(n6863), .A2(n5189), .Y(n6906) );
  NAND2X0_RVT U6245 ( .A1(n6864), .A2(n4960), .Y(n6904) );
  NAND3X0_RVT U6246 ( .A1(n6907), .A2(n6908), .A3(n6909), .Y(n4684) );
  NAND2X0_RVT U6247 ( .A1(n6863), .A2(n5174), .Y(n6909) );
  NAND2X0_RVT U6248 ( .A1(n6910), .A2(Datai[15]), .Y(n6908) );
  NAND2X0_RVT U6249 ( .A1(n6864), .A2(n4945), .Y(n6907) );
  NAND4X0_RVT U6250 ( .A1(n6911), .A2(n6912), .A3(n6913), .A4(n6914), .Y(n4683) );
  NAND2X0_RVT U6251 ( .A1(n5203), .A2(n5088), .Y(n6914) );
  NAND2X0_RVT U6252 ( .A1(n6915), .A2(n5211), .Y(n6913) );
  NAND2X0_RVT U6253 ( .A1(n5196), .A2(Datai[16]), .Y(n6912) );
  NAND2X0_RVT U6254 ( .A1(n6916), .A2(n5210), .Y(n6911) );
  NAND4X0_RVT U6255 ( .A1(n6917), .A2(n6918), .A3(n6919), .A4(n6920), .Y(n4682) );
  NAND2X0_RVT U6256 ( .A1(n5202), .A2(n5087), .Y(n6920) );
  NAND2X0_RVT U6257 ( .A1(n6921), .A2(n5209), .Y(n6919) );
  NAND2X0_RVT U6258 ( .A1(n5199), .A2(Datai[17]), .Y(n6918) );
  NAND2X0_RVT U6259 ( .A1(n6922), .A2(n5208), .Y(n6917) );
  NAND4X0_RVT U6260 ( .A1(n6923), .A2(n6924), .A3(n6925), .A4(n6926), .Y(n4681) );
  NAND2X0_RVT U6261 ( .A1(n5201), .A2(n5089), .Y(n6926) );
  NAND2X0_RVT U6262 ( .A1(n6927), .A2(n5211), .Y(n6925) );
  NAND2X0_RVT U6263 ( .A1(n5198), .A2(Datai[18]), .Y(n6924) );
  NAND2X0_RVT U6264 ( .A1(n6928), .A2(n5210), .Y(n6923) );
  NAND4X0_RVT U6265 ( .A1(n6929), .A2(n6930), .A3(n6931), .A4(n6932), .Y(n4680) );
  NAND2X0_RVT U6266 ( .A1(n5200), .A2(n5090), .Y(n6932) );
  NAND2X0_RVT U6267 ( .A1(n6933), .A2(n5209), .Y(n6931) );
  NAND2X0_RVT U6268 ( .A1(n5197), .A2(Datai[19]), .Y(n6930) );
  NAND2X0_RVT U6269 ( .A1(n6934), .A2(n5208), .Y(n6929) );
  NAND4X0_RVT U6270 ( .A1(n6935), .A2(n6936), .A3(n6937), .A4(n6938), .Y(n4679) );
  NAND2X0_RVT U6271 ( .A1(n5203), .A2(n5091), .Y(n6938) );
  NAND2X0_RVT U6272 ( .A1(n6939), .A2(n5211), .Y(n6937) );
  NAND2X0_RVT U6273 ( .A1(n5196), .A2(Datai[20]), .Y(n6936) );
  NAND2X0_RVT U6274 ( .A1(n6940), .A2(n5210), .Y(n6935) );
  NAND4X0_RVT U6275 ( .A1(n6941), .A2(n6942), .A3(n6943), .A4(n6944), .Y(n4678) );
  NAND2X0_RVT U6276 ( .A1(n5202), .A2(n5092), .Y(n6944) );
  NAND2X0_RVT U6277 ( .A1(n6945), .A2(n5209), .Y(n6943) );
  NAND2X0_RVT U6278 ( .A1(n5199), .A2(Datai[21]), .Y(n6942) );
  NAND2X0_RVT U6279 ( .A1(n6946), .A2(n5208), .Y(n6941) );
  NAND4X0_RVT U6280 ( .A1(n6947), .A2(n6948), .A3(n6949), .A4(n6950), .Y(n4677) );
  NAND2X0_RVT U6281 ( .A1(n5201), .A2(n5093), .Y(n6950) );
  NAND2X0_RVT U6282 ( .A1(n6951), .A2(n5211), .Y(n6949) );
  NAND2X0_RVT U6283 ( .A1(n5198), .A2(Datai[22]), .Y(n6948) );
  NAND2X0_RVT U6284 ( .A1(n6952), .A2(n5210), .Y(n6947) );
  NAND4X0_RVT U6285 ( .A1(n6953), .A2(n6954), .A3(n6955), .A4(n6956), .Y(n4676) );
  NAND2X0_RVT U6286 ( .A1(n5200), .A2(n5094), .Y(n6956) );
  NAND2X0_RVT U6287 ( .A1(n6957), .A2(n5209), .Y(n6955) );
  NAND2X0_RVT U6288 ( .A1(n5197), .A2(Datai[23]), .Y(n6954) );
  NAND2X0_RVT U6289 ( .A1(n6958), .A2(n5208), .Y(n6953) );
  NAND4X0_RVT U6290 ( .A1(n6959), .A2(n6960), .A3(n6961), .A4(n6962), .Y(n4675) );
  NAND2X0_RVT U6291 ( .A1(n5203), .A2(n5095), .Y(n6962) );
  NAND2X0_RVT U6292 ( .A1(n6963), .A2(n5211), .Y(n6961) );
  NAND2X0_RVT U6293 ( .A1(n5196), .A2(Datai[24]), .Y(n6960) );
  NAND2X0_RVT U6294 ( .A1(n6964), .A2(n5210), .Y(n6959) );
  NAND4X0_RVT U6295 ( .A1(n6965), .A2(n6966), .A3(n6967), .A4(n6968), .Y(n4674) );
  NAND2X0_RVT U6296 ( .A1(n5202), .A2(n5096), .Y(n6968) );
  NAND2X0_RVT U6297 ( .A1(n6969), .A2(n5209), .Y(n6967) );
  NAND2X0_RVT U6298 ( .A1(Datai[25]), .A2(n5199), .Y(n6966) );
  NAND2X0_RVT U6299 ( .A1(n6970), .A2(n5208), .Y(n6965) );
  NAND4X0_RVT U6300 ( .A1(n6971), .A2(n6972), .A3(n6973), .A4(n6974), .Y(n4673) );
  NAND2X0_RVT U6301 ( .A1(n5201), .A2(n5097), .Y(n6974) );
  NAND2X0_RVT U6302 ( .A1(n6975), .A2(n5211), .Y(n6973) );
  NAND2X0_RVT U6303 ( .A1(Datai[26]), .A2(n5198), .Y(n6972) );
  NAND2X0_RVT U6304 ( .A1(n6976), .A2(n5210), .Y(n6971) );
  NAND4X0_RVT U6305 ( .A1(n6977), .A2(n6978), .A3(n6979), .A4(n6980), .Y(n4672) );
  NAND2X0_RVT U6306 ( .A1(n5200), .A2(n5098), .Y(n6980) );
  NAND2X0_RVT U6307 ( .A1(n6981), .A2(n5209), .Y(n6979) );
  NAND2X0_RVT U6308 ( .A1(Datai[27]), .A2(n5197), .Y(n6978) );
  NAND2X0_RVT U6309 ( .A1(n6982), .A2(n5208), .Y(n6977) );
  NAND4X0_RVT U6310 ( .A1(n6983), .A2(n6984), .A3(n6985), .A4(n6986), .Y(n4671) );
  NAND2X0_RVT U6311 ( .A1(n5203), .A2(n5099), .Y(n6986) );
  NAND2X0_RVT U6312 ( .A1(n6987), .A2(n5211), .Y(n6985) );
  NAND2X0_RVT U6313 ( .A1(n5199), .A2(Datai[28]), .Y(n6984) );
  NAND2X0_RVT U6314 ( .A1(n6988), .A2(n5210), .Y(n6983) );
  NAND4X0_RVT U6315 ( .A1(n6989), .A2(n6990), .A3(n6991), .A4(n6992), .Y(n4670) );
  NAND2X0_RVT U6316 ( .A1(n5202), .A2(n5100), .Y(n6992) );
  NAND2X0_RVT U6317 ( .A1(n6993), .A2(n5209), .Y(n6991) );
  NAND2X0_RVT U6318 ( .A1(n5198), .A2(Datai[29]), .Y(n6990) );
  NAND2X0_RVT U6319 ( .A1(n6994), .A2(n5208), .Y(n6989) );
  NAND4X0_RVT U6320 ( .A1(n6995), .A2(n6996), .A3(n6997), .A4(n6998), .Y(n4669) );
  NAND2X0_RVT U6321 ( .A1(n5201), .A2(n5101), .Y(n6998) );
  NAND2X0_RVT U6322 ( .A1(n6999), .A2(n5211), .Y(n6997) );
  NAND2X0_RVT U6323 ( .A1(n5197), .A2(Datai[30]), .Y(n6996) );
  NAND2X0_RVT U6324 ( .A1(n7000), .A2(n5210), .Y(n6995) );
  NAND3X0_RVT U6325 ( .A1(n7001), .A2(n7002), .A3(n7003), .Y(n4668) );
  NAND2X0_RVT U6326 ( .A1(n5200), .A2(n5054), .Y(n7003) );
  NAND2X0_RVT U6327 ( .A1(n5196), .A2(Datai[31]), .Y(n7002) );
  NAND4X0_RVT U6328 ( .A1(n7005), .A2(n7006), .A3(n7007), .A4(n7008), .Y(n6768) );
  NAND3X0_RVT U6329 ( .A1(n7009), .A2(n5268), .A3(n7004), .Y(n7005) );
  INVX0_RVT U6330 ( .A(n7010), .Y(n7004) );
  XNOR2X1_RVT U6331 ( .A1(n7011), .A2(n7012), .Y(n7001) );
  NAND2X0_RVT U6332 ( .A1(n7013), .A2(n7014), .Y(n7012) );
  NAND2X0_RVT U6333 ( .A1(n5207), .A2(n5054), .Y(n7011) );
  NAND3X0_RVT U6334 ( .A1(n7015), .A2(n6861), .A3(n7016), .Y(n4667) );
  NAND2X0_RVT U6335 ( .A1(uWord[0]), .A2(n6863), .Y(n7016) );
  NAND2X0_RVT U6336 ( .A1(n6910), .A2(Datai[0]), .Y(n6861) );
  NAND2X0_RVT U6337 ( .A1(n6864), .A2(n6769), .Y(n7015) );
  NAND3X0_RVT U6338 ( .A1(n7017), .A2(n6866), .A3(n7018), .Y(n4666) );
  NAND2X0_RVT U6339 ( .A1(uWord[1]), .A2(n6863), .Y(n7018) );
  NAND2X0_RVT U6340 ( .A1(n6910), .A2(Datai[1]), .Y(n6866) );
  NAND2X0_RVT U6341 ( .A1(n6864), .A2(n6775), .Y(n7017) );
  NAND3X0_RVT U6342 ( .A1(n7019), .A2(n6869), .A3(n7020), .Y(n4665) );
  NAND2X0_RVT U6343 ( .A1(uWord[2]), .A2(n6863), .Y(n7020) );
  NAND2X0_RVT U6344 ( .A1(n6910), .A2(Datai[2]), .Y(n6869) );
  NAND2X0_RVT U6345 ( .A1(n6864), .A2(n6781), .Y(n7019) );
  NAND3X0_RVT U6346 ( .A1(n7021), .A2(n6872), .A3(n7022), .Y(n4664) );
  NAND2X0_RVT U6347 ( .A1(uWord[3]), .A2(n6863), .Y(n7022) );
  NAND2X0_RVT U6348 ( .A1(n6910), .A2(Datai[3]), .Y(n6872) );
  NAND2X0_RVT U6349 ( .A1(n6864), .A2(n6787), .Y(n7021) );
  NAND3X0_RVT U6350 ( .A1(n7023), .A2(n6875), .A3(n7024), .Y(n4663) );
  NAND2X0_RVT U6351 ( .A1(uWord[4]), .A2(n6863), .Y(n7024) );
  NAND2X0_RVT U6352 ( .A1(n6910), .A2(Datai[4]), .Y(n6875) );
  NAND2X0_RVT U6353 ( .A1(n6864), .A2(n6793), .Y(n7023) );
  NAND3X0_RVT U6354 ( .A1(n7025), .A2(n6878), .A3(n7026), .Y(n4662) );
  NAND2X0_RVT U6355 ( .A1(uWord[5]), .A2(n6863), .Y(n7026) );
  NAND2X0_RVT U6356 ( .A1(n6910), .A2(Datai[5]), .Y(n6878) );
  NAND2X0_RVT U6357 ( .A1(n6864), .A2(n6799), .Y(n7025) );
  NAND3X0_RVT U6358 ( .A1(n7027), .A2(n6881), .A3(n7028), .Y(n4661) );
  NAND2X0_RVT U6359 ( .A1(uWord[6]), .A2(n6863), .Y(n7028) );
  NAND2X0_RVT U6360 ( .A1(n6910), .A2(Datai[6]), .Y(n6881) );
  NAND2X0_RVT U6361 ( .A1(n6864), .A2(n6805), .Y(n7027) );
  NAND3X0_RVT U6362 ( .A1(n7029), .A2(n6884), .A3(n7030), .Y(n4660) );
  NAND2X0_RVT U6363 ( .A1(uWord[7]), .A2(n6863), .Y(n7030) );
  NAND2X0_RVT U6364 ( .A1(n6910), .A2(Datai[7]), .Y(n6884) );
  NAND2X0_RVT U6365 ( .A1(n6864), .A2(n6811), .Y(n7029) );
  NAND3X0_RVT U6366 ( .A1(n7031), .A2(n6887), .A3(n7032), .Y(n4659) );
  NAND2X0_RVT U6367 ( .A1(uWord[8]), .A2(n6863), .Y(n7032) );
  NAND2X0_RVT U6368 ( .A1(n6910), .A2(Datai[8]), .Y(n6887) );
  NAND2X0_RVT U6369 ( .A1(n6864), .A2(n6817), .Y(n7031) );
  NAND3X0_RVT U6370 ( .A1(n7033), .A2(n6890), .A3(n7034), .Y(n4658) );
  NAND2X0_RVT U6371 ( .A1(uWord[9]), .A2(n6863), .Y(n7034) );
  NAND2X0_RVT U6372 ( .A1(n6910), .A2(Datai[9]), .Y(n6890) );
  NAND2X0_RVT U6373 ( .A1(n6864), .A2(n6823), .Y(n7033) );
  NAND3X0_RVT U6374 ( .A1(n7035), .A2(n6893), .A3(n7036), .Y(n4657) );
  NAND2X0_RVT U6375 ( .A1(uWord[10]), .A2(n6863), .Y(n7036) );
  NAND2X0_RVT U6376 ( .A1(n6910), .A2(Datai[10]), .Y(n6893) );
  NAND2X0_RVT U6377 ( .A1(n6864), .A2(n6829), .Y(n7035) );
  NAND3X0_RVT U6378 ( .A1(n7037), .A2(n6896), .A3(n7038), .Y(n4656) );
  NAND2X0_RVT U6379 ( .A1(uWord[11]), .A2(n6863), .Y(n7038) );
  NAND2X0_RVT U6380 ( .A1(n6910), .A2(Datai[11]), .Y(n6896) );
  NAND2X0_RVT U6381 ( .A1(n6864), .A2(n6835), .Y(n7037) );
  NAND3X0_RVT U6382 ( .A1(n7039), .A2(n6899), .A3(n7040), .Y(n4655) );
  NAND2X0_RVT U6383 ( .A1(uWord[12]), .A2(n6863), .Y(n7040) );
  NAND2X0_RVT U6384 ( .A1(n6910), .A2(Datai[12]), .Y(n6899) );
  NAND2X0_RVT U6385 ( .A1(n6864), .A2(n6841), .Y(n7039) );
  NAND3X0_RVT U6386 ( .A1(n7041), .A2(n6902), .A3(n7042), .Y(n4654) );
  NAND2X0_RVT U6387 ( .A1(uWord[13]), .A2(n6863), .Y(n7042) );
  NAND2X0_RVT U6388 ( .A1(n6910), .A2(Datai[13]), .Y(n6902) );
  NAND2X0_RVT U6389 ( .A1(n6864), .A2(n6847), .Y(n7041) );
  NAND3X0_RVT U6390 ( .A1(n7043), .A2(n6905), .A3(n7044), .Y(n4653) );
  NAND2X0_RVT U6391 ( .A1(uWord[14]), .A2(n6863), .Y(n7044) );
  NAND2X0_RVT U6392 ( .A1(n6910), .A2(Datai[14]), .Y(n6905) );
  AND2X1_RVT U6393 ( .A1(n7046), .A2(n7045), .Y(n6910) );
  NAND2X0_RVT U6394 ( .A1(n6864), .A2(n6853), .Y(n7043) );
  NAND2X0_RVT U6395 ( .A1(n7047), .A2(n7008), .Y(n7045) );
  NAND3X0_RVT U6396 ( .A1(n7048), .A2(n7049), .A3(n7050), .Y(n4652) );
  NAND2X0_RVT U6397 ( .A1(n7051), .A2(n4911), .Y(n7049) );
  NAND2X0_RVT U6398 ( .A1(n6767), .A2(n7052), .Y(n7048) );
  NAND3X0_RVT U6399 ( .A1(n7053), .A2(n7054), .A3(n7055), .Y(n4651) );
  NAND2X0_RVT U6400 ( .A1(n6774), .A2(n7052), .Y(n7055) );
  NAND2X0_RVT U6401 ( .A1(n7056), .A2(n4964), .Y(n7054) );
  NAND2X0_RVT U6402 ( .A1(n7052), .A2(n7050), .Y(n7056) );
  NAND2X0_RVT U6403 ( .A1(n9544), .A2(n7057), .Y(n7050) );
  NAND3X0_RVT U6404 ( .A1(n7057), .A2(n4911), .A3(n9543), .Y(n7053) );
  NAND3X0_RVT U6405 ( .A1(n7058), .A2(n7059), .A3(n7060), .Y(n4650) );
  NAND2X0_RVT U6406 ( .A1(n7057), .A2(n7061), .Y(n7060) );
  XNOR2X1_RVT U6407 ( .A1(n7062), .A2(n4940), .Y(n7061) );
  NAND2X0_RVT U6408 ( .A1(n7051), .A2(n4940), .Y(n7059) );
  NAND2X0_RVT U6409 ( .A1(n6780), .A2(n7052), .Y(n7058) );
  NAND3X0_RVT U6410 ( .A1(n7063), .A2(n7064), .A3(n7065), .Y(n4649) );
  NAND2X0_RVT U6411 ( .A1(n7057), .A2(n7066), .Y(n7065) );
  XNOR2X1_RVT U6412 ( .A1(n7067), .A2(n4939), .Y(n7066) );
  NAND2X0_RVT U6413 ( .A1(n7051), .A2(n4939), .Y(n7064) );
  NAND2X0_RVT U6414 ( .A1(n6786), .A2(n7052), .Y(n7063) );
  NAND3X0_RVT U6415 ( .A1(n7068), .A2(n7069), .A3(n7070), .Y(n4648) );
  NAND2X0_RVT U6416 ( .A1(n7057), .A2(n7071), .Y(n7070) );
  XNOR2X1_RVT U6417 ( .A1(n7072), .A2(n4941), .Y(n7071) );
  NAND2X0_RVT U6418 ( .A1(n7051), .A2(n4941), .Y(n7069) );
  NAND2X0_RVT U6419 ( .A1(n6792), .A2(n7052), .Y(n7068) );
  NAND3X0_RVT U6420 ( .A1(n7073), .A2(n7074), .A3(n7075), .Y(n4647) );
  NAND2X0_RVT U6421 ( .A1(n7057), .A2(n7076), .Y(n7075) );
  XNOR2X1_RVT U6422 ( .A1(n7077), .A2(n4938), .Y(n7076) );
  NAND2X0_RVT U6423 ( .A1(n7051), .A2(n4938), .Y(n7074) );
  NAND2X0_RVT U6424 ( .A1(n6798), .A2(n7052), .Y(n7073) );
  NAND3X0_RVT U6425 ( .A1(n7078), .A2(n7079), .A3(n7080), .Y(n4646) );
  NAND2X0_RVT U6426 ( .A1(n7057), .A2(n7081), .Y(n7080) );
  XNOR2X1_RVT U6427 ( .A1(n7082), .A2(n4942), .Y(n7081) );
  NAND2X0_RVT U6428 ( .A1(n7051), .A2(n4942), .Y(n7079) );
  NAND2X0_RVT U6429 ( .A1(n6804), .A2(n7052), .Y(n7078) );
  NAND3X0_RVT U6430 ( .A1(n7083), .A2(n7084), .A3(n7085), .Y(n4645) );
  NAND2X0_RVT U6431 ( .A1(n7057), .A2(n7086), .Y(n7085) );
  XNOR2X1_RVT U6432 ( .A1(n7087), .A2(n4937), .Y(n7086) );
  NAND2X0_RVT U6433 ( .A1(n7051), .A2(n4937), .Y(n7084) );
  NAND2X0_RVT U6434 ( .A1(n6810), .A2(n7052), .Y(n7083) );
  NAND3X0_RVT U6435 ( .A1(n7088), .A2(n7089), .A3(n7090), .Y(n4644) );
  NAND2X0_RVT U6436 ( .A1(n7057), .A2(n7091), .Y(n7090) );
  XNOR2X1_RVT U6437 ( .A1(n7092), .A2(n4943), .Y(n7091) );
  NAND2X0_RVT U6438 ( .A1(n7051), .A2(n4943), .Y(n7089) );
  NAND2X0_RVT U6439 ( .A1(n6816), .A2(n7052), .Y(n7088) );
  NAND3X0_RVT U6440 ( .A1(n7093), .A2(n7094), .A3(n7095), .Y(n4643) );
  NAND2X0_RVT U6441 ( .A1(n7057), .A2(n7096), .Y(n7095) );
  XNOR2X1_RVT U6442 ( .A1(n7097), .A2(n4933), .Y(n7096) );
  NAND2X0_RVT U6443 ( .A1(n7051), .A2(n4933), .Y(n7094) );
  NAND2X0_RVT U6444 ( .A1(n6822), .A2(n7052), .Y(n7093) );
  NAND3X0_RVT U6445 ( .A1(n7098), .A2(n7099), .A3(n7100), .Y(n4642) );
  NAND2X0_RVT U6446 ( .A1(n7057), .A2(n7101), .Y(n7100) );
  XOR2X1_RVT U6447 ( .A1(n7102), .A2(n7103), .Y(n7101) );
  NAND2X0_RVT U6448 ( .A1(n7051), .A2(n4966), .Y(n7099) );
  NAND2X0_RVT U6449 ( .A1(n6828), .A2(n7052), .Y(n7098) );
  NAND3X0_RVT U6450 ( .A1(n7104), .A2(n7105), .A3(n7106), .Y(n4641) );
  NAND2X0_RVT U6451 ( .A1(n7057), .A2(n7107), .Y(n7106) );
  XNOR2X1_RVT U6452 ( .A1(n7108), .A2(n4936), .Y(n7107) );
  NAND2X0_RVT U6453 ( .A1(n7051), .A2(n4936), .Y(n7105) );
  NAND2X0_RVT U6454 ( .A1(n6834), .A2(n7052), .Y(n7104) );
  NAND3X0_RVT U6455 ( .A1(n7109), .A2(n7110), .A3(n7111), .Y(n4640) );
  NAND2X0_RVT U6456 ( .A1(n7057), .A2(n7112), .Y(n7111) );
  XNOR2X1_RVT U6457 ( .A1(n7113), .A2(n4944), .Y(n7112) );
  NAND2X0_RVT U6458 ( .A1(n7051), .A2(n4944), .Y(n7110) );
  NAND2X0_RVT U6459 ( .A1(n6840), .A2(n7052), .Y(n7109) );
  NAND3X0_RVT U6460 ( .A1(n7114), .A2(n7115), .A3(n7116), .Y(n4639) );
  NAND2X0_RVT U6461 ( .A1(n7057), .A2(n7117), .Y(n7116) );
  XNOR2X1_RVT U6462 ( .A1(n7118), .A2(n4935), .Y(n7117) );
  NAND2X0_RVT U6463 ( .A1(n7051), .A2(n4935), .Y(n7115) );
  NAND2X0_RVT U6464 ( .A1(n6846), .A2(n7052), .Y(n7114) );
  NAND3X0_RVT U6465 ( .A1(n7119), .A2(n7120), .A3(n7121), .Y(n4638) );
  NAND2X0_RVT U6466 ( .A1(n7057), .A2(n7122), .Y(n7121) );
  XNOR2X1_RVT U6467 ( .A1(n7123), .A2(n4934), .Y(n7122) );
  NAND2X0_RVT U6468 ( .A1(n7051), .A2(n4934), .Y(n7120) );
  NAND2X0_RVT U6469 ( .A1(n6852), .A2(n7052), .Y(n7119) );
  NAND3X0_RVT U6470 ( .A1(n7124), .A2(n7125), .A3(n7126), .Y(n4637) );
  NAND2X0_RVT U6471 ( .A1(n7057), .A2(n7127), .Y(n7126) );
  XNOR2X1_RVT U6472 ( .A1(n7128), .A2(n4932), .Y(n7127) );
  NAND2X0_RVT U6473 ( .A1(n7051), .A2(n4932), .Y(n7125) );
  NAND2X0_RVT U6474 ( .A1(n6858), .A2(n7052), .Y(n7124) );
  NAND3X0_RVT U6475 ( .A1(n7129), .A2(n7130), .A3(n7131), .Y(n4636) );
  NAND2X0_RVT U6476 ( .A1(n7057), .A2(n7132), .Y(n7131) );
  NAND2X0_RVT U6477 ( .A1(n7051), .A2(n4986), .Y(n7130) );
  NAND2X0_RVT U6478 ( .A1(n6915), .A2(n7052), .Y(n7129) );
  NAND3X0_RVT U6479 ( .A1(n7133), .A2(n7134), .A3(n7135), .Y(n4635) );
  NAND2X0_RVT U6480 ( .A1(n7057), .A2(n7136), .Y(n7135) );
  NAND2X0_RVT U6481 ( .A1(n7051), .A2(n4987), .Y(n7134) );
  NAND2X0_RVT U6482 ( .A1(n6921), .A2(n7052), .Y(n7133) );
  NAND3X0_RVT U6483 ( .A1(n7137), .A2(n7138), .A3(n7139), .Y(n4634) );
  NAND2X0_RVT U6484 ( .A1(n7057), .A2(n7140), .Y(n7139) );
  NAND2X0_RVT U6485 ( .A1(n7051), .A2(n4992), .Y(n7138) );
  NAND2X0_RVT U6486 ( .A1(n6927), .A2(n7052), .Y(n7137) );
  NAND3X0_RVT U6487 ( .A1(n7141), .A2(n7142), .A3(n7143), .Y(n4633) );
  NAND2X0_RVT U6488 ( .A1(n7057), .A2(n7144), .Y(n7143) );
  NAND2X0_RVT U6489 ( .A1(n7051), .A2(n4993), .Y(n7142) );
  NAND2X0_RVT U6490 ( .A1(n6933), .A2(n7052), .Y(n7141) );
  NAND3X0_RVT U6491 ( .A1(n7145), .A2(n7146), .A3(n7147), .Y(n4632) );
  NAND2X0_RVT U6492 ( .A1(n7057), .A2(n7148), .Y(n7147) );
  NAND2X0_RVT U6493 ( .A1(n7051), .A2(n4994), .Y(n7146) );
  NAND2X0_RVT U6494 ( .A1(n6939), .A2(n7052), .Y(n7145) );
  NAND3X0_RVT U6495 ( .A1(n7149), .A2(n7150), .A3(n7151), .Y(n4631) );
  NAND2X0_RVT U6496 ( .A1(n7057), .A2(n7152), .Y(n7151) );
  NAND2X0_RVT U6497 ( .A1(n7051), .A2(n4995), .Y(n7150) );
  NAND2X0_RVT U6498 ( .A1(n6945), .A2(n7052), .Y(n7149) );
  NAND3X0_RVT U6499 ( .A1(n7153), .A2(n7154), .A3(n7155), .Y(n4630) );
  NAND2X0_RVT U6500 ( .A1(n7057), .A2(n7156), .Y(n7155) );
  NAND2X0_RVT U6501 ( .A1(n7051), .A2(n4991), .Y(n7154) );
  NAND2X0_RVT U6502 ( .A1(n6951), .A2(n7052), .Y(n7153) );
  NAND3X0_RVT U6503 ( .A1(n7157), .A2(n7158), .A3(n7159), .Y(n4629) );
  NAND2X0_RVT U6504 ( .A1(n7057), .A2(n7160), .Y(n7159) );
  NAND2X0_RVT U6505 ( .A1(n7051), .A2(n4990), .Y(n7158) );
  NAND2X0_RVT U6506 ( .A1(n6957), .A2(n7052), .Y(n7157) );
  NAND3X0_RVT U6507 ( .A1(n7161), .A2(n7162), .A3(n7163), .Y(n4628) );
  NAND2X0_RVT U6508 ( .A1(n7057), .A2(n7164), .Y(n7163) );
  NAND2X0_RVT U6509 ( .A1(n7051), .A2(n4985), .Y(n7162) );
  NAND2X0_RVT U6510 ( .A1(n6963), .A2(n7052), .Y(n7161) );
  NAND3X0_RVT U6511 ( .A1(n7165), .A2(n7166), .A3(n7167), .Y(n4627) );
  NAND2X0_RVT U6512 ( .A1(n7057), .A2(n7168), .Y(n7167) );
  NAND2X0_RVT U6513 ( .A1(n7051), .A2(n4984), .Y(n7166) );
  NAND2X0_RVT U6514 ( .A1(n6969), .A2(n7052), .Y(n7165) );
  NAND3X0_RVT U6515 ( .A1(n7169), .A2(n7170), .A3(n7171), .Y(n4626) );
  NAND2X0_RVT U6516 ( .A1(n7057), .A2(n7172), .Y(n7171) );
  NAND2X0_RVT U6517 ( .A1(n7051), .A2(n4983), .Y(n7170) );
  NAND2X0_RVT U6518 ( .A1(n6975), .A2(n7052), .Y(n7169) );
  NAND3X0_RVT U6519 ( .A1(n7173), .A2(n7174), .A3(n7175), .Y(n4625) );
  NAND2X0_RVT U6520 ( .A1(n7057), .A2(n7176), .Y(n7175) );
  NAND2X0_RVT U6521 ( .A1(n7051), .A2(n4982), .Y(n7174) );
  NAND2X0_RVT U6522 ( .A1(n6981), .A2(n7052), .Y(n7173) );
  NAND3X0_RVT U6523 ( .A1(n7177), .A2(n7178), .A3(n7179), .Y(n4624) );
  NAND2X0_RVT U6524 ( .A1(n7057), .A2(n7180), .Y(n7179) );
  NAND2X0_RVT U6525 ( .A1(n7051), .A2(n4981), .Y(n7178) );
  NAND2X0_RVT U6526 ( .A1(n6987), .A2(n7052), .Y(n7177) );
  NAND3X0_RVT U6527 ( .A1(n7181), .A2(n7182), .A3(n7183), .Y(n4623) );
  NAND2X0_RVT U6528 ( .A1(n7057), .A2(n7184), .Y(n7183) );
  NAND2X0_RVT U6529 ( .A1(n7051), .A2(n4980), .Y(n7182) );
  NAND2X0_RVT U6530 ( .A1(n6993), .A2(n7052), .Y(n7181) );
  NAND3X0_RVT U6531 ( .A1(n7185), .A2(n7186), .A3(n7187), .Y(n4622) );
  NAND2X0_RVT U6532 ( .A1(n7057), .A2(n7188), .Y(n7187) );
  NAND2X0_RVT U6533 ( .A1(n7051), .A2(n4988), .Y(n7186) );
  NAND2X0_RVT U6534 ( .A1(n6999), .A2(n7052), .Y(n7185) );
  NAND2X0_RVT U6535 ( .A1(n7189), .A2(n7190), .Y(n4621) );
  NAND2X0_RVT U6536 ( .A1(n7191), .A2(n7057), .Y(n7190) );
  XNOR2X1_RVT U6537 ( .A1(n7193), .A2(n4958), .Y(n7191) );
  NAND2X0_RVT U6538 ( .A1(n7194), .A2(n7195), .Y(n7193) );
  INVX0_RVT U6539 ( .A(n7196), .Y(n7194) );
  NAND2X0_RVT U6540 ( .A1(n7051), .A2(n4958), .Y(n7189) );
  NAND2X0_RVT U6541 ( .A1(n7192), .A2(n5265), .Y(n7198) );
  NAND4X0_RVT U6542 ( .A1(n7199), .A2(n7200), .A3(n7201), .A4(n7202), .Y(n4620) );
  AND4X1_RVT U6543 ( .A1(n7203), .A2(n7204), .A3(n7205), .A4(n7206), .Y(n7202)
         );
  NAND2X0_RVT U6544 ( .A1(n7207), .A2(n5397), .Y(n7206) );
  XOR2X1_RVT U6545 ( .A1(n7208), .A2(n7209), .Y(n5397) );
  NAND2X0_RVT U6546 ( .A1(n7210), .A2(n7211), .Y(n7205) );
  NAND2X0_RVT U6547 ( .A1(n7212), .A2(n4911), .Y(n7204) );
  NAND2X0_RVT U6548 ( .A1(n7213), .A2(n7214), .Y(n7203) );
  NAND2X0_RVT U6549 ( .A1(n7215), .A2(n5055), .Y(n7201) );
  NAND2X0_RVT U6550 ( .A1(n6767), .A2(n5371), .Y(n7200) );
  XNOR2X1_RVT U6551 ( .A1(n7216), .A2(n7217), .Y(n6767) );
  NAND2X0_RVT U6552 ( .A1(n7218), .A2(rEIP[0]), .Y(n7199) );
  NAND4X0_RVT U6553 ( .A1(n7219), .A2(n7220), .A3(n7221), .A4(n7222), .Y(n4619) );
  AND4X1_RVT U6554 ( .A1(n7223), .A2(n7224), .A3(n7225), .A4(n7226), .Y(n7222)
         );
  NAND2X0_RVT U6555 ( .A1(n7207), .A2(n5411), .Y(n7226) );
  XOR2X1_RVT U6556 ( .A1(n7227), .A2(n7228), .Y(n5411) );
  NAND2X0_RVT U6557 ( .A1(n7229), .A2(n7230), .Y(n7227) );
  NAND2X0_RVT U6558 ( .A1(n7212), .A2(n4964), .Y(n7225) );
  NAND2X0_RVT U6559 ( .A1(n7231), .A2(n7210), .Y(n7224) );
  NAND2X0_RVT U6560 ( .A1(n7232), .A2(n7214), .Y(n7223) );
  NAND2X0_RVT U6561 ( .A1(n7215), .A2(n5063), .Y(n7221) );
  NAND2X0_RVT U6562 ( .A1(n5371), .A2(n6774), .Y(n7220) );
  XOR2X1_RVT U6563 ( .A1(n7233), .A2(n7234), .Y(n6774) );
  NAND2X0_RVT U6564 ( .A1(n7218), .A2(rEIP[1]), .Y(n7219) );
  NAND4X0_RVT U6565 ( .A1(n7235), .A2(n7236), .A3(n7237), .A4(n7238), .Y(n4618) );
  AND4X1_RVT U6566 ( .A1(n7239), .A2(n7240), .A3(n7241), .A4(n7242), .Y(n7238)
         );
  NAND2X0_RVT U6567 ( .A1(n7207), .A2(n5421), .Y(n7242) );
  XNOR2X1_RVT U6568 ( .A1(n7243), .A2(n7244), .Y(n5421) );
  NAND2X0_RVT U6569 ( .A1(n7245), .A2(n7246), .Y(n7243) );
  NAND2X0_RVT U6570 ( .A1(n7247), .A2(n7210), .Y(n7241) );
  NAND2X0_RVT U6571 ( .A1(n7212), .A2(n4940), .Y(n7240) );
  NAND2X0_RVT U6572 ( .A1(n7248), .A2(n7214), .Y(n7239) );
  NAND2X0_RVT U6573 ( .A1(n7215), .A2(n5062), .Y(n7237) );
  NAND2X0_RVT U6574 ( .A1(n5371), .A2(n6780), .Y(n7236) );
  XOR2X1_RVT U6575 ( .A1(n7249), .A2(n7250), .Y(n6780) );
  NAND2X0_RVT U6576 ( .A1(n7218), .A2(rEIP[2]), .Y(n7235) );
  NAND4X0_RVT U6577 ( .A1(n7251), .A2(n7252), .A3(n7253), .A4(n7254), .Y(n4617) );
  AND4X1_RVT U6578 ( .A1(n7255), .A2(n7256), .A3(n7257), .A4(n7258), .Y(n7254)
         );
  NAND2X0_RVT U6579 ( .A1(n7207), .A2(n5431), .Y(n7258) );
  NAND2X0_RVT U6580 ( .A1(n7260), .A2(n7261), .Y(n6377) );
  OR2X1_RVT U6581 ( .A1(n7246), .A2(n7244), .Y(n7261) );
  NAND2X0_RVT U6582 ( .A1(n7262), .A2(n4926), .Y(n7246) );
  OR2X1_RVT U6583 ( .A1(n7245), .A2(n7244), .Y(n7260) );
  AND2X1_RVT U6584 ( .A1(n7263), .A2(n7264), .Y(n7244) );
  NAND2X0_RVT U6585 ( .A1(n7265), .A2(n7228), .Y(n7264) );
  INVX0_RVT U6586 ( .A(n7230), .Y(n7265) );
  NAND2X0_RVT U6587 ( .A1(n7262), .A2(n4927), .Y(n7230) );
  NAND2X0_RVT U6588 ( .A1(n7266), .A2(n7228), .Y(n7263) );
  AND2X1_RVT U6589 ( .A1(n7208), .A2(n7209), .Y(n7228) );
  NAND3X0_RVT U6590 ( .A1(n7267), .A2(n7268), .A3(n7269), .Y(n7209) );
  NAND2X0_RVT U6591 ( .A1(n7262), .A2(n4908), .Y(n7269) );
  NAND2X0_RVT U6592 ( .A1(n6310), .A2(n6529), .Y(n7268) );
  OR2X1_RVT U6593 ( .A1(n7270), .A2(n7271), .Y(n6529) );
  OR4X1_RVT U6594 ( .A1(Datai[0]), .A2(Datai[1]), .A3(Datai[2]), .A4(Datai[3]), 
        .Y(n7271) );
  OR4X1_RVT U6595 ( .A1(Datai[4]), .A2(Datai[5]), .A3(Datai[6]), .A4(Datai[7]), 
        .Y(n7270) );
  AND2X1_RVT U6596 ( .A1(Datai[31]), .A2(n5476), .Y(n6310) );
  OR2X1_RVT U6597 ( .A1(n6523), .A2(n5390), .Y(n7267) );
  NAND2X0_RVT U6598 ( .A1(Datai[31]), .A2(n7272), .Y(n6523) );
  OR2X1_RVT U6599 ( .A1(n7273), .A2(n7274), .Y(n7272) );
  OR4X1_RVT U6600 ( .A1(Datai[10]), .A2(Datai[11]), .A3(Datai[12]), .A4(
        Datai[13]), .Y(n7274) );
  OR4X1_RVT U6601 ( .A1(Datai[14]), .A2(Datai[15]), .A3(Datai[8]), .A4(
        Datai[9]), .Y(n7273) );
  NAND2X0_RVT U6602 ( .A1(n7275), .A2(n7276), .Y(n7208) );
  NAND2X0_RVT U6603 ( .A1(Datai[16]), .A2(n5476), .Y(n7276) );
  INVX0_RVT U6604 ( .A(n7262), .Y(n7275) );
  INVX0_RVT U6605 ( .A(n7229), .Y(n7266) );
  NAND2X0_RVT U6606 ( .A1(Datai[17]), .A2(n5476), .Y(n7229) );
  NAND2X0_RVT U6607 ( .A1(Datai[18]), .A2(n5476), .Y(n7245) );
  NAND2X0_RVT U6608 ( .A1(n6378), .A2(n7277), .Y(n7259) );
  NAND2X0_RVT U6609 ( .A1(n7262), .A2(n4906), .Y(n7277) );
  NAND2X0_RVT U6610 ( .A1(n7278), .A2(n5363), .Y(n7262) );
  NAND2X0_RVT U6611 ( .A1(n6306), .A2(n6434), .Y(n5363) );
  NAND2X0_RVT U6612 ( .A1(n7009), .A2(n7279), .Y(n7278) );
  NAND2X0_RVT U6613 ( .A1(Datai[19]), .A2(n5476), .Y(n6378) );
  NAND2X0_RVT U6614 ( .A1(n7212), .A2(n4939), .Y(n7257) );
  NAND2X0_RVT U6615 ( .A1(n7280), .A2(n7210), .Y(n7256) );
  NAND2X0_RVT U6616 ( .A1(n7281), .A2(n7214), .Y(n7255) );
  NAND2X0_RVT U6617 ( .A1(n7215), .A2(n5061), .Y(n7253) );
  NAND2X0_RVT U6618 ( .A1(n5371), .A2(n6786), .Y(n7252) );
  XOR2X1_RVT U6619 ( .A1(n7282), .A2(n7283), .Y(n6786) );
  NAND2X0_RVT U6620 ( .A1(n7218), .A2(rEIP[3]), .Y(n7251) );
  NAND4X0_RVT U6621 ( .A1(n7284), .A2(n7285), .A3(n7286), .A4(n7287), .Y(n4616) );
  AND4X1_RVT U6622 ( .A1(n7288), .A2(n7289), .A3(n7290), .A4(n6433), .Y(n7287)
         );
  NAND2X0_RVT U6623 ( .A1(n7291), .A2(n7210), .Y(n7290) );
  NAND2X0_RVT U6624 ( .A1(n7212), .A2(n4941), .Y(n7289) );
  NAND2X0_RVT U6625 ( .A1(n7292), .A2(n7214), .Y(n7288) );
  NAND2X0_RVT U6626 ( .A1(n7215), .A2(n5060), .Y(n7286) );
  NAND2X0_RVT U6627 ( .A1(n5371), .A2(n6792), .Y(n7285) );
  XOR2X1_RVT U6628 ( .A1(n7293), .A2(n7294), .Y(n6792) );
  NAND2X0_RVT U6629 ( .A1(n7218), .A2(rEIP[4]), .Y(n7284) );
  NAND4X0_RVT U6630 ( .A1(n7295), .A2(n7296), .A3(n7297), .A4(n7298), .Y(n4615) );
  AND4X1_RVT U6631 ( .A1(n7299), .A2(n7300), .A3(n7301), .A4(n6433), .Y(n7298)
         );
  NAND2X0_RVT U6632 ( .A1(n7212), .A2(n4938), .Y(n7301) );
  NAND2X0_RVT U6633 ( .A1(n7302), .A2(n7210), .Y(n7300) );
  NAND2X0_RVT U6634 ( .A1(n7303), .A2(n7214), .Y(n7299) );
  NAND2X0_RVT U6635 ( .A1(n7215), .A2(n5059), .Y(n7297) );
  NAND2X0_RVT U6636 ( .A1(n5371), .A2(n6798), .Y(n7296) );
  XOR2X1_RVT U6637 ( .A1(n7304), .A2(n7305), .Y(n6798) );
  NAND2X0_RVT U6638 ( .A1(n7218), .A2(rEIP[5]), .Y(n7295) );
  NAND4X0_RVT U6639 ( .A1(n7306), .A2(n7307), .A3(n7308), .A4(n7309), .Y(n4614) );
  AND4X1_RVT U6640 ( .A1(n7310), .A2(n7311), .A3(n7312), .A4(n6433), .Y(n7309)
         );
  NAND2X0_RVT U6641 ( .A1(n7313), .A2(n7210), .Y(n7312) );
  NAND2X0_RVT U6642 ( .A1(n7212), .A2(n4942), .Y(n7311) );
  NAND2X0_RVT U6643 ( .A1(n7314), .A2(n7214), .Y(n7310) );
  NAND2X0_RVT U6644 ( .A1(n7215), .A2(n5058), .Y(n7308) );
  NAND2X0_RVT U6645 ( .A1(n5371), .A2(n6804), .Y(n7307) );
  XOR2X1_RVT U6646 ( .A1(n7315), .A2(n7316), .Y(n6804) );
  NAND2X0_RVT U6647 ( .A1(n7218), .A2(rEIP[6]), .Y(n7306) );
  NAND4X0_RVT U6648 ( .A1(n7317), .A2(n7318), .A3(n7319), .A4(n7320), .Y(n4613) );
  AND4X1_RVT U6649 ( .A1(n7321), .A2(n7322), .A3(n7323), .A4(n6433), .Y(n7320)
         );
  NAND2X0_RVT U6650 ( .A1(n7212), .A2(n4937), .Y(n7323) );
  NAND2X0_RVT U6651 ( .A1(n7324), .A2(n7210), .Y(n7322) );
  NAND2X0_RVT U6652 ( .A1(n7325), .A2(n7214), .Y(n7321) );
  NAND2X0_RVT U6653 ( .A1(n7215), .A2(n5057), .Y(n7319) );
  NAND2X0_RVT U6654 ( .A1(n5371), .A2(n6810), .Y(n7318) );
  XOR2X1_RVT U6655 ( .A1(n7326), .A2(n7327), .Y(n6810) );
  NAND2X0_RVT U6656 ( .A1(n7218), .A2(rEIP[7]), .Y(n7317) );
  NAND4X0_RVT U6657 ( .A1(n7328), .A2(n7329), .A3(n7330), .A4(n7331), .Y(n4612) );
  AND4X1_RVT U6658 ( .A1(n7332), .A2(n7333), .A3(n7334), .A4(n6433), .Y(n7331)
         );
  NAND2X0_RVT U6659 ( .A1(n7335), .A2(n7210), .Y(n7334) );
  NAND2X0_RVT U6660 ( .A1(n7212), .A2(n4943), .Y(n7333) );
  NAND2X0_RVT U6661 ( .A1(n7336), .A2(n7214), .Y(n7332) );
  NAND2X0_RVT U6662 ( .A1(n7215), .A2(n5064), .Y(n7330) );
  NAND2X0_RVT U6663 ( .A1(n5371), .A2(n6816), .Y(n7329) );
  XOR2X1_RVT U6664 ( .A1(n7337), .A2(n7338), .Y(n6816) );
  NAND2X0_RVT U6665 ( .A1(n7218), .A2(rEIP[8]), .Y(n7328) );
  NAND4X0_RVT U6666 ( .A1(n7339), .A2(n7340), .A3(n7341), .A4(n7342), .Y(n4611) );
  AND4X1_RVT U6667 ( .A1(n7343), .A2(n7344), .A3(n7345), .A4(n6433), .Y(n7342)
         );
  NAND2X0_RVT U6668 ( .A1(n7212), .A2(n4933), .Y(n7345) );
  NAND2X0_RVT U6669 ( .A1(n7346), .A2(n7210), .Y(n7344) );
  NAND2X0_RVT U6670 ( .A1(n7347), .A2(n7214), .Y(n7343) );
  NAND2X0_RVT U6671 ( .A1(n7215), .A2(n5065), .Y(n7341) );
  NAND2X0_RVT U6672 ( .A1(n5371), .A2(n6822), .Y(n7340) );
  XOR2X1_RVT U6673 ( .A1(n7348), .A2(n7349), .Y(n6822) );
  NAND2X0_RVT U6674 ( .A1(n7218), .A2(rEIP[9]), .Y(n7339) );
  NAND4X0_RVT U6675 ( .A1(n7350), .A2(n7351), .A3(n7352), .A4(n7353), .Y(n4610) );
  AND4X1_RVT U6676 ( .A1(n7354), .A2(n7355), .A3(n7356), .A4(n6433), .Y(n7353)
         );
  NAND2X0_RVT U6677 ( .A1(n7357), .A2(n7210), .Y(n7356) );
  NAND2X0_RVT U6678 ( .A1(n7212), .A2(n4966), .Y(n7355) );
  NAND2X0_RVT U6679 ( .A1(n7358), .A2(n7214), .Y(n7354) );
  NAND2X0_RVT U6680 ( .A1(n7215), .A2(n5066), .Y(n7352) );
  NAND2X0_RVT U6681 ( .A1(n5371), .A2(n6828), .Y(n7351) );
  XOR2X1_RVT U6682 ( .A1(n7359), .A2(n7360), .Y(n6828) );
  NAND2X0_RVT U6683 ( .A1(n7218), .A2(rEIP[10]), .Y(n7350) );
  NAND4X0_RVT U6684 ( .A1(n7361), .A2(n7362), .A3(n7363), .A4(n7364), .Y(n4609) );
  AND4X1_RVT U6685 ( .A1(n7365), .A2(n7366), .A3(n7367), .A4(n6433), .Y(n7364)
         );
  NAND2X0_RVT U6686 ( .A1(n7212), .A2(n4936), .Y(n7367) );
  NAND2X0_RVT U6687 ( .A1(n7368), .A2(n7210), .Y(n7366) );
  NAND2X0_RVT U6688 ( .A1(n7369), .A2(n7214), .Y(n7365) );
  NAND2X0_RVT U6689 ( .A1(n7215), .A2(n5067), .Y(n7363) );
  NAND2X0_RVT U6690 ( .A1(n5371), .A2(n6834), .Y(n7362) );
  XOR2X1_RVT U6691 ( .A1(n7370), .A2(n7371), .Y(n6834) );
  NAND2X0_RVT U6692 ( .A1(n7218), .A2(rEIP[11]), .Y(n7361) );
  NAND4X0_RVT U6693 ( .A1(n7372), .A2(n7373), .A3(n7374), .A4(n7375), .Y(n4608) );
  AND4X1_RVT U6694 ( .A1(n7376), .A2(n7377), .A3(n7378), .A4(n6433), .Y(n7375)
         );
  NAND2X0_RVT U6695 ( .A1(n7379), .A2(n7210), .Y(n7378) );
  NAND2X0_RVT U6696 ( .A1(n7212), .A2(n4944), .Y(n7377) );
  NAND2X0_RVT U6697 ( .A1(n7380), .A2(n7214), .Y(n7376) );
  NAND2X0_RVT U6698 ( .A1(n7215), .A2(n5068), .Y(n7374) );
  NAND2X0_RVT U6699 ( .A1(n5371), .A2(n6840), .Y(n7373) );
  XOR2X1_RVT U6700 ( .A1(n7381), .A2(n7382), .Y(n6840) );
  NAND2X0_RVT U6701 ( .A1(n7218), .A2(rEIP[12]), .Y(n7372) );
  NAND4X0_RVT U6702 ( .A1(n7383), .A2(n7384), .A3(n7385), .A4(n7386), .Y(n4607) );
  AND4X1_RVT U6703 ( .A1(n7387), .A2(n7388), .A3(n7389), .A4(n6433), .Y(n7386)
         );
  NAND2X0_RVT U6704 ( .A1(n7212), .A2(n4935), .Y(n7389) );
  NAND2X0_RVT U6705 ( .A1(n7390), .A2(n7210), .Y(n7388) );
  NAND2X0_RVT U6706 ( .A1(n7391), .A2(n7214), .Y(n7387) );
  NAND2X0_RVT U6707 ( .A1(n7215), .A2(n5069), .Y(n7385) );
  NAND2X0_RVT U6708 ( .A1(n5371), .A2(n6846), .Y(n7384) );
  XOR2X1_RVT U6709 ( .A1(n7392), .A2(n7393), .Y(n6846) );
  NAND2X0_RVT U6710 ( .A1(n7218), .A2(rEIP[13]), .Y(n7383) );
  NAND4X0_RVT U6711 ( .A1(n7394), .A2(n7395), .A3(n7396), .A4(n7397), .Y(n4606) );
  AND4X1_RVT U6712 ( .A1(n7398), .A2(n7399), .A3(n7400), .A4(n6433), .Y(n7397)
         );
  NAND2X0_RVT U6713 ( .A1(n7401), .A2(n7210), .Y(n7400) );
  NAND2X0_RVT U6714 ( .A1(n7212), .A2(n4934), .Y(n7399) );
  NAND2X0_RVT U6715 ( .A1(n7402), .A2(n7214), .Y(n7398) );
  NAND2X0_RVT U6716 ( .A1(n7215), .A2(n5070), .Y(n7396) );
  NAND2X0_RVT U6717 ( .A1(n5371), .A2(n6852), .Y(n7395) );
  XOR2X1_RVT U6718 ( .A1(n7403), .A2(n7404), .Y(n6852) );
  NAND2X0_RVT U6719 ( .A1(n7218), .A2(rEIP[14]), .Y(n7394) );
  NAND4X0_RVT U6720 ( .A1(n7405), .A2(n7406), .A3(n7407), .A4(n7408), .Y(n4605) );
  AND4X1_RVT U6721 ( .A1(n7409), .A2(n7410), .A3(n7411), .A4(n6433), .Y(n7408)
         );
  NAND2X0_RVT U6722 ( .A1(n7212), .A2(n4932), .Y(n7411) );
  NAND2X0_RVT U6723 ( .A1(n7412), .A2(n7210), .Y(n7410) );
  NAND2X0_RVT U6724 ( .A1(n7413), .A2(n7214), .Y(n7409) );
  NAND2X0_RVT U6725 ( .A1(n7215), .A2(n5071), .Y(n7407) );
  NAND2X0_RVT U6726 ( .A1(n5371), .A2(n6858), .Y(n7406) );
  XOR2X1_RVT U6727 ( .A1(n7414), .A2(n7415), .Y(n6858) );
  NAND2X0_RVT U6728 ( .A1(n7218), .A2(rEIP[15]), .Y(n7405) );
  NAND4X0_RVT U6729 ( .A1(n7416), .A2(n7417), .A3(n7418), .A4(n7419), .Y(n4604) );
  AND4X1_RVT U6730 ( .A1(n7420), .A2(n7421), .A3(n7422), .A4(n6433), .Y(n7419)
         );
  NAND2X0_RVT U6731 ( .A1(n7212), .A2(n4986), .Y(n7422) );
  NAND2X0_RVT U6732 ( .A1(n7210), .A2(n7423), .Y(n7421) );
  NAND2X0_RVT U6733 ( .A1(n7424), .A2(n7214), .Y(n7420) );
  NAND2X0_RVT U6734 ( .A1(n7215), .A2(n5072), .Y(n7418) );
  NAND2X0_RVT U6735 ( .A1(n5371), .A2(n6915), .Y(n7417) );
  NAND3X0_RVT U6736 ( .A1(n7425), .A2(n7426), .A3(n7427), .Y(n6915) );
  XNOR2X1_RVT U6737 ( .A1(n7428), .A2(n7429), .Y(n7427) );
  NAND2X0_RVT U6738 ( .A1(n7132), .A2(n7430), .Y(n7426) );
  XOR2X1_RVT U6739 ( .A1(n7431), .A2(n7432), .Y(n7132) );
  NAND2X0_RVT U6740 ( .A1(n7218), .A2(rEIP[16]), .Y(n7416) );
  NAND4X0_RVT U6741 ( .A1(n7433), .A2(n7434), .A3(n7435), .A4(n7436), .Y(n4603) );
  AND4X1_RVT U6742 ( .A1(n7437), .A2(n7438), .A3(n7439), .A4(n6433), .Y(n7436)
         );
  NAND2X0_RVT U6743 ( .A1(n7212), .A2(n4987), .Y(n7439) );
  NAND2X0_RVT U6744 ( .A1(n7440), .A2(n7210), .Y(n7438) );
  NAND2X0_RVT U6745 ( .A1(n7441), .A2(n7214), .Y(n7437) );
  NAND2X0_RVT U6746 ( .A1(n7215), .A2(n5073), .Y(n7435) );
  NAND2X0_RVT U6747 ( .A1(n5371), .A2(n6921), .Y(n7434) );
  NAND3X0_RVT U6748 ( .A1(n7442), .A2(n7443), .A3(n7444), .Y(n6921) );
  XNOR2X1_RVT U6749 ( .A1(n7445), .A2(n7446), .Y(n7444) );
  NAND2X0_RVT U6750 ( .A1(n7136), .A2(n7430), .Y(n7443) );
  XNOR2X1_RVT U6751 ( .A1(n7447), .A2(n7448), .Y(n7136) );
  NAND2X0_RVT U6752 ( .A1(n7431), .A2(n7432), .Y(n7447) );
  NAND2X0_RVT U6753 ( .A1(n7218), .A2(rEIP[17]), .Y(n7433) );
  NAND4X0_RVT U6754 ( .A1(n7449), .A2(n7450), .A3(n7451), .A4(n7452), .Y(n4602) );
  AND4X1_RVT U6755 ( .A1(n7453), .A2(n7454), .A3(n7455), .A4(n6433), .Y(n7452)
         );
  NAND2X0_RVT U6756 ( .A1(n7212), .A2(n4992), .Y(n7455) );
  NAND2X0_RVT U6757 ( .A1(n7456), .A2(n7210), .Y(n7454) );
  NAND2X0_RVT U6758 ( .A1(n7457), .A2(n7214), .Y(n7453) );
  NAND2X0_RVT U6759 ( .A1(n7215), .A2(n5074), .Y(n7451) );
  NAND2X0_RVT U6760 ( .A1(n5371), .A2(n6927), .Y(n7450) );
  NAND3X0_RVT U6761 ( .A1(n7458), .A2(n7459), .A3(n7460), .Y(n6927) );
  XNOR2X1_RVT U6762 ( .A1(n7461), .A2(n7462), .Y(n7460) );
  NAND2X0_RVT U6763 ( .A1(n7140), .A2(n7430), .Y(n7459) );
  XOR2X1_RVT U6764 ( .A1(n7463), .A2(n7464), .Y(n7140) );
  NAND2X0_RVT U6765 ( .A1(n7218), .A2(rEIP[18]), .Y(n7449) );
  NAND4X0_RVT U6766 ( .A1(n7465), .A2(n7466), .A3(n7467), .A4(n7468), .Y(n4601) );
  AND4X1_RVT U6767 ( .A1(n7469), .A2(n7470), .A3(n7471), .A4(n6433), .Y(n7468)
         );
  NAND2X0_RVT U6768 ( .A1(n7212), .A2(n4993), .Y(n7471) );
  NAND2X0_RVT U6769 ( .A1(n7472), .A2(n7210), .Y(n7470) );
  NAND2X0_RVT U6770 ( .A1(n7473), .A2(n7214), .Y(n7469) );
  NAND2X0_RVT U6771 ( .A1(n7215), .A2(n5075), .Y(n7467) );
  NAND2X0_RVT U6772 ( .A1(n5371), .A2(n6933), .Y(n7466) );
  NAND3X0_RVT U6773 ( .A1(n7474), .A2(n7475), .A3(n7476), .Y(n6933) );
  XNOR2X1_RVT U6774 ( .A1(n7477), .A2(n7478), .Y(n7476) );
  NAND2X0_RVT U6775 ( .A1(n7144), .A2(n7430), .Y(n7475) );
  XNOR2X1_RVT U6776 ( .A1(n7479), .A2(n7480), .Y(n7144) );
  NAND2X0_RVT U6777 ( .A1(n7463), .A2(n7464), .Y(n7479) );
  NAND2X0_RVT U6778 ( .A1(n7218), .A2(rEIP[19]), .Y(n7465) );
  NAND4X0_RVT U6779 ( .A1(n7481), .A2(n7482), .A3(n7483), .A4(n7484), .Y(n4600) );
  AND3X1_RVT U6780 ( .A1(n7485), .A2(n7486), .A3(n7487), .Y(n7484) );
  NAND2X0_RVT U6781 ( .A1(n7488), .A2(n7214), .Y(n7487) );
  NAND2X0_RVT U6782 ( .A1(n7212), .A2(n4994), .Y(n7486) );
  NAND2X0_RVT U6783 ( .A1(n7489), .A2(n7210), .Y(n7485) );
  NAND2X0_RVT U6784 ( .A1(n7215), .A2(n5076), .Y(n7483) );
  NAND2X0_RVT U6785 ( .A1(n5371), .A2(n6939), .Y(n7482) );
  NAND3X0_RVT U6786 ( .A1(n7490), .A2(n7491), .A3(n7492), .Y(n6939) );
  XNOR2X1_RVT U6787 ( .A1(n7493), .A2(n7494), .Y(n7492) );
  NAND2X0_RVT U6788 ( .A1(n7148), .A2(n7430), .Y(n7491) );
  XOR2X1_RVT U6789 ( .A1(n7495), .A2(n7496), .Y(n7148) );
  NAND2X0_RVT U6790 ( .A1(n7218), .A2(rEIP[20]), .Y(n7481) );
  NAND4X0_RVT U6791 ( .A1(n7497), .A2(n7498), .A3(n7499), .A4(n7500), .Y(n4599) );
  AND3X1_RVT U6792 ( .A1(n7501), .A2(n7502), .A3(n7503), .Y(n7500) );
  NAND2X0_RVT U6793 ( .A1(n7504), .A2(n7214), .Y(n7503) );
  NAND2X0_RVT U6794 ( .A1(n7212), .A2(n4995), .Y(n7502) );
  NAND2X0_RVT U6795 ( .A1(n7505), .A2(n7210), .Y(n7501) );
  NAND2X0_RVT U6796 ( .A1(n7215), .A2(n5077), .Y(n7499) );
  NAND2X0_RVT U6797 ( .A1(n5371), .A2(n6945), .Y(n7498) );
  NAND3X0_RVT U6798 ( .A1(n7506), .A2(n7507), .A3(n7508), .Y(n6945) );
  XNOR2X1_RVT U6799 ( .A1(n7509), .A2(n7510), .Y(n7508) );
  NAND2X0_RVT U6800 ( .A1(n7152), .A2(n7430), .Y(n7507) );
  XNOR2X1_RVT U6801 ( .A1(n7511), .A2(n7512), .Y(n7152) );
  NAND2X0_RVT U6802 ( .A1(n7495), .A2(n7496), .Y(n7511) );
  NAND2X0_RVT U6803 ( .A1(n7218), .A2(rEIP[21]), .Y(n7497) );
  NAND4X0_RVT U6804 ( .A1(n7513), .A2(n7514), .A3(n7515), .A4(n7516), .Y(n4598) );
  AND3X1_RVT U6805 ( .A1(n7517), .A2(n7518), .A3(n7519), .Y(n7516) );
  NAND2X0_RVT U6806 ( .A1(n7520), .A2(n7214), .Y(n7519) );
  NAND2X0_RVT U6807 ( .A1(n7212), .A2(n4991), .Y(n7518) );
  NAND2X0_RVT U6808 ( .A1(n7521), .A2(n7210), .Y(n7517) );
  NAND2X0_RVT U6809 ( .A1(n7215), .A2(n5078), .Y(n7515) );
  NAND2X0_RVT U6810 ( .A1(n5371), .A2(n6951), .Y(n7514) );
  NAND3X0_RVT U6811 ( .A1(n7522), .A2(n7523), .A3(n7524), .Y(n6951) );
  XNOR2X1_RVT U6812 ( .A1(n7525), .A2(n7526), .Y(n7524) );
  NAND2X0_RVT U6813 ( .A1(n7156), .A2(n7430), .Y(n7523) );
  XOR2X1_RVT U6814 ( .A1(n7527), .A2(n7528), .Y(n7156) );
  NAND2X0_RVT U6815 ( .A1(n7218), .A2(rEIP[22]), .Y(n7513) );
  NAND4X0_RVT U6816 ( .A1(n7529), .A2(n7530), .A3(n7531), .A4(n7532), .Y(n4597) );
  AND3X1_RVT U6817 ( .A1(n7533), .A2(n7534), .A3(n7535), .Y(n7532) );
  NAND2X0_RVT U6818 ( .A1(n7536), .A2(n7214), .Y(n7535) );
  NAND2X0_RVT U6819 ( .A1(n7212), .A2(n4990), .Y(n7534) );
  NAND2X0_RVT U6820 ( .A1(n7537), .A2(n7210), .Y(n7533) );
  NAND2X0_RVT U6821 ( .A1(n7215), .A2(n5079), .Y(n7531) );
  NAND2X0_RVT U6822 ( .A1(n5371), .A2(n6957), .Y(n7530) );
  NAND3X0_RVT U6823 ( .A1(n7538), .A2(n7539), .A3(n7540), .Y(n6957) );
  XNOR2X1_RVT U6824 ( .A1(n7541), .A2(n7542), .Y(n7540) );
  NAND2X0_RVT U6825 ( .A1(n7160), .A2(n7430), .Y(n7539) );
  XOR3X1_RVT U6826 ( .A1(n7543), .A2(n7544), .A3(n7545), .Y(n7160) );
  NAND2X0_RVT U6827 ( .A1(n7218), .A2(rEIP[23]), .Y(n7529) );
  NAND4X0_RVT U6828 ( .A1(n7546), .A2(n7547), .A3(n7548), .A4(n7549), .Y(n4596) );
  AND3X1_RVT U6829 ( .A1(n7550), .A2(n7551), .A3(n7552), .Y(n7549) );
  NAND2X0_RVT U6830 ( .A1(n7553), .A2(n7214), .Y(n7552) );
  NAND2X0_RVT U6831 ( .A1(n7212), .A2(n4985), .Y(n7551) );
  NAND2X0_RVT U6832 ( .A1(n7554), .A2(n7210), .Y(n7550) );
  NAND2X0_RVT U6833 ( .A1(n7215), .A2(n5080), .Y(n7548) );
  NAND2X0_RVT U6834 ( .A1(n5371), .A2(n6963), .Y(n7547) );
  NAND3X0_RVT U6835 ( .A1(n7555), .A2(n7556), .A3(n7557), .Y(n6963) );
  XNOR2X1_RVT U6836 ( .A1(n7558), .A2(n7559), .Y(n7557) );
  NAND2X0_RVT U6837 ( .A1(n7164), .A2(n7430), .Y(n7556) );
  XOR2X1_RVT U6838 ( .A1(n7560), .A2(n7561), .Y(n7164) );
  OR2X1_RVT U6839 ( .A1(n7562), .A2(n7563), .Y(n7560) );
  NAND2X0_RVT U6840 ( .A1(n7218), .A2(rEIP[24]), .Y(n7546) );
  NAND4X0_RVT U6841 ( .A1(n7564), .A2(n7565), .A3(n7566), .A4(n7567), .Y(n4595) );
  AND3X1_RVT U6842 ( .A1(n7568), .A2(n7569), .A3(n7570), .Y(n7567) );
  NAND2X0_RVT U6843 ( .A1(n7571), .A2(n7214), .Y(n7570) );
  NAND2X0_RVT U6844 ( .A1(n7212), .A2(n4984), .Y(n7569) );
  NAND2X0_RVT U6845 ( .A1(n7572), .A2(n7210), .Y(n7568) );
  NAND2X0_RVT U6846 ( .A1(n7215), .A2(n5081), .Y(n7566) );
  NAND2X0_RVT U6847 ( .A1(n5371), .A2(n6969), .Y(n7565) );
  NAND3X0_RVT U6848 ( .A1(n7573), .A2(n7574), .A3(n7575), .Y(n6969) );
  XNOR2X1_RVT U6849 ( .A1(n7576), .A2(n7577), .Y(n7575) );
  NAND2X0_RVT U6850 ( .A1(n7168), .A2(n7430), .Y(n7574) );
  XOR2X1_RVT U6851 ( .A1(n7578), .A2(n7579), .Y(n7168) );
  OR2X1_RVT U6852 ( .A1(n7580), .A2(n7581), .Y(n7578) );
  NAND2X0_RVT U6853 ( .A1(n7218), .A2(rEIP[25]), .Y(n7564) );
  NAND4X0_RVT U6854 ( .A1(n7582), .A2(n7583), .A3(n7584), .A4(n7585), .Y(n4594) );
  AND3X1_RVT U6855 ( .A1(n7586), .A2(n7587), .A3(n7588), .Y(n7585) );
  NAND2X0_RVT U6856 ( .A1(n7589), .A2(n7214), .Y(n7588) );
  NAND2X0_RVT U6857 ( .A1(n7212), .A2(n4983), .Y(n7587) );
  NAND2X0_RVT U6858 ( .A1(n7590), .A2(n7210), .Y(n7586) );
  NAND2X0_RVT U6859 ( .A1(n7215), .A2(n5082), .Y(n7584) );
  NAND2X0_RVT U6860 ( .A1(n5371), .A2(n6975), .Y(n7583) );
  NAND3X0_RVT U6861 ( .A1(n7591), .A2(n7592), .A3(n7593), .Y(n6975) );
  XNOR2X1_RVT U6862 ( .A1(n7594), .A2(n7595), .Y(n7593) );
  NAND2X0_RVT U6863 ( .A1(n7172), .A2(n7430), .Y(n7592) );
  XOR2X1_RVT U6864 ( .A1(n7596), .A2(n7597), .Y(n7172) );
  OR2X1_RVT U6865 ( .A1(n7598), .A2(n7599), .Y(n7596) );
  NAND2X0_RVT U6866 ( .A1(n7218), .A2(rEIP[26]), .Y(n7582) );
  NAND4X0_RVT U6867 ( .A1(n7600), .A2(n7601), .A3(n7602), .A4(n7603), .Y(n4593) );
  AND3X1_RVT U6868 ( .A1(n7604), .A2(n7605), .A3(n7606), .Y(n7603) );
  NAND2X0_RVT U6869 ( .A1(n7607), .A2(n7214), .Y(n7606) );
  NAND2X0_RVT U6870 ( .A1(n7212), .A2(n4982), .Y(n7605) );
  NAND2X0_RVT U6871 ( .A1(n7608), .A2(n7210), .Y(n7604) );
  NAND2X0_RVT U6872 ( .A1(n7215), .A2(n5083), .Y(n7602) );
  NAND2X0_RVT U6873 ( .A1(n5371), .A2(n6981), .Y(n7601) );
  NAND3X0_RVT U6874 ( .A1(n7609), .A2(n7610), .A3(n7611), .Y(n6981) );
  XNOR2X1_RVT U6875 ( .A1(n7612), .A2(n7613), .Y(n7611) );
  NAND2X0_RVT U6876 ( .A1(n7176), .A2(n7430), .Y(n7610) );
  XOR2X1_RVT U6877 ( .A1(n7614), .A2(n7615), .Y(n7176) );
  OR2X1_RVT U6878 ( .A1(n7616), .A2(n7617), .Y(n7614) );
  NAND2X0_RVT U6879 ( .A1(n7218), .A2(rEIP[27]), .Y(n7600) );
  NAND4X0_RVT U6880 ( .A1(n7618), .A2(n7619), .A3(n7620), .A4(n7621), .Y(n4592) );
  AND3X1_RVT U6881 ( .A1(n7622), .A2(n7623), .A3(n7624), .Y(n7621) );
  NAND2X0_RVT U6882 ( .A1(n7625), .A2(n7214), .Y(n7624) );
  NAND2X0_RVT U6883 ( .A1(n7212), .A2(n4981), .Y(n7623) );
  NAND2X0_RVT U6884 ( .A1(n7626), .A2(n7210), .Y(n7622) );
  NAND2X0_RVT U6885 ( .A1(n7215), .A2(n5084), .Y(n7620) );
  NAND2X0_RVT U6886 ( .A1(n5371), .A2(n6987), .Y(n7619) );
  NAND3X0_RVT U6887 ( .A1(n7627), .A2(n7628), .A3(n7629), .Y(n6987) );
  XNOR2X1_RVT U6888 ( .A1(n7630), .A2(n7631), .Y(n7629) );
  NAND2X0_RVT U6889 ( .A1(n7180), .A2(n7430), .Y(n7628) );
  XOR2X1_RVT U6890 ( .A1(n7632), .A2(n7633), .Y(n7180) );
  OR2X1_RVT U6891 ( .A1(n7634), .A2(n7635), .Y(n7632) );
  NAND2X0_RVT U6892 ( .A1(n7218), .A2(rEIP[28]), .Y(n7618) );
  NAND4X0_RVT U6893 ( .A1(n7636), .A2(n7637), .A3(n7638), .A4(n7639), .Y(n4591) );
  AND3X1_RVT U6894 ( .A1(n7640), .A2(n7641), .A3(n7642), .Y(n7639) );
  NAND2X0_RVT U6895 ( .A1(n7643), .A2(n7214), .Y(n7642) );
  NAND2X0_RVT U6896 ( .A1(n7212), .A2(n4980), .Y(n7641) );
  NAND2X0_RVT U6897 ( .A1(n7644), .A2(n7210), .Y(n7640) );
  NAND2X0_RVT U6898 ( .A1(n7215), .A2(n5085), .Y(n7638) );
  NAND2X0_RVT U6899 ( .A1(n5371), .A2(n6993), .Y(n7637) );
  NAND3X0_RVT U6900 ( .A1(n7645), .A2(n7646), .A3(n7647), .Y(n6993) );
  XNOR2X1_RVT U6901 ( .A1(n7648), .A2(n7649), .Y(n7647) );
  NAND2X0_RVT U6902 ( .A1(n7184), .A2(n7430), .Y(n7646) );
  XOR2X1_RVT U6903 ( .A1(n7650), .A2(n7651), .Y(n7184) );
  OR2X1_RVT U6904 ( .A1(n7652), .A2(n7653), .Y(n7650) );
  NAND2X0_RVT U6905 ( .A1(n7218), .A2(rEIP[29]), .Y(n7636) );
  NAND4X0_RVT U6906 ( .A1(n7654), .A2(n7655), .A3(n7656), .A4(n7657), .Y(n4590) );
  AND3X1_RVT U6907 ( .A1(n7658), .A2(n7659), .A3(n7660), .Y(n7657) );
  NAND2X0_RVT U6908 ( .A1(n7661), .A2(n7214), .Y(n7660) );
  NAND2X0_RVT U6909 ( .A1(n7212), .A2(n4988), .Y(n7659) );
  NAND2X0_RVT U6910 ( .A1(n7662), .A2(n7210), .Y(n7658) );
  NAND2X0_RVT U6911 ( .A1(n7215), .A2(n5056), .Y(n7656) );
  NAND2X0_RVT U6912 ( .A1(n5371), .A2(n6999), .Y(n7655) );
  NAND3X0_RVT U6913 ( .A1(n7663), .A2(n7664), .A3(n7665), .Y(n6999) );
  XNOR2X1_RVT U6914 ( .A1(n7666), .A2(n7667), .Y(n7665) );
  NAND2X0_RVT U6915 ( .A1(n7188), .A2(n7430), .Y(n7664) );
  XOR2X1_RVT U6916 ( .A1(n7668), .A2(n7195), .Y(n7188) );
  NAND2X0_RVT U6917 ( .A1(n7669), .A2(n7670), .Y(n7195) );
  NAND2X0_RVT U6918 ( .A1(n7653), .A2(n7651), .Y(n7670) );
  AND2X1_RVT U6919 ( .A1(n7192), .A2(n4980), .Y(n7653) );
  NAND2X0_RVT U6920 ( .A1(n7651), .A2(n7652), .Y(n7669) );
  NAND4X0_RVT U6921 ( .A1(n7671), .A2(n7672), .A3(n7673), .A4(n7674), .Y(n7652) );
  NAND2X0_RVT U6922 ( .A1(n7675), .A2(n7676), .Y(n7674) );
  NAND2X0_RVT U6923 ( .A1(n873), .A2(n7677), .Y(n7676) );
  NAND2X0_RVT U6924 ( .A1(n7678), .A2(n5042), .Y(n7677) );
  NAND2X0_RVT U6925 ( .A1(n7679), .A2(n7680), .Y(n7673) );
  NAND2X0_RVT U6926 ( .A1(n7681), .A2(n7682), .Y(n7672) );
  NAND2X0_RVT U6927 ( .A1(n7683), .A2(n7684), .Y(n7671) );
  NAND2X0_RVT U6928 ( .A1(n7685), .A2(n7686), .Y(n7651) );
  NAND2X0_RVT U6929 ( .A1(n7635), .A2(n7633), .Y(n7686) );
  AND2X1_RVT U6930 ( .A1(n7192), .A2(n4981), .Y(n7635) );
  NAND2X0_RVT U6931 ( .A1(n7633), .A2(n7634), .Y(n7685) );
  NAND4X0_RVT U6932 ( .A1(n7687), .A2(n7688), .A3(n7689), .A4(n7690), .Y(n7634) );
  NAND2X0_RVT U6933 ( .A1(n7675), .A2(n7691), .Y(n7690) );
  NAND2X0_RVT U6934 ( .A1(n7692), .A2(n7693), .Y(n7691) );
  NAND2X0_RVT U6935 ( .A1(n7694), .A2(n5036), .Y(n7693) );
  NAND2X0_RVT U6936 ( .A1(n7678), .A2(n5035), .Y(n7692) );
  NAND2X0_RVT U6937 ( .A1(n7679), .A2(n7695), .Y(n7689) );
  NAND2X0_RVT U6938 ( .A1(n7681), .A2(n7696), .Y(n7688) );
  NAND2X0_RVT U6939 ( .A1(n7683), .A2(n7697), .Y(n7687) );
  NAND2X0_RVT U6940 ( .A1(n7698), .A2(n7699), .Y(n7633) );
  NAND2X0_RVT U6941 ( .A1(n7617), .A2(n7615), .Y(n7699) );
  AND2X1_RVT U6942 ( .A1(n7192), .A2(n4982), .Y(n7617) );
  NAND2X0_RVT U6943 ( .A1(n7615), .A2(n7616), .Y(n7698) );
  NAND4X0_RVT U6944 ( .A1(n7700), .A2(n7701), .A3(n7702), .A4(n7703), .Y(n7616) );
  NAND2X0_RVT U6945 ( .A1(n7675), .A2(n7704), .Y(n7703) );
  NAND2X0_RVT U6946 ( .A1(n7705), .A2(n7706), .Y(n7704) );
  NAND2X0_RVT U6947 ( .A1(n7694), .A2(n5029), .Y(n7706) );
  NAND2X0_RVT U6948 ( .A1(n7678), .A2(n5028), .Y(n7705) );
  NAND2X0_RVT U6949 ( .A1(n7679), .A2(n7707), .Y(n7702) );
  NAND2X0_RVT U6950 ( .A1(n7681), .A2(n7708), .Y(n7701) );
  NAND2X0_RVT U6951 ( .A1(n7683), .A2(n7709), .Y(n7700) );
  NAND2X0_RVT U6952 ( .A1(n7710), .A2(n7711), .Y(n7615) );
  NAND2X0_RVT U6953 ( .A1(n7599), .A2(n7597), .Y(n7711) );
  AND2X1_RVT U6954 ( .A1(n7192), .A2(n4983), .Y(n7599) );
  NAND2X0_RVT U6955 ( .A1(n7597), .A2(n7598), .Y(n7710) );
  NAND4X0_RVT U6956 ( .A1(n7712), .A2(n7713), .A3(n7714), .A4(n7715), .Y(n7598) );
  NAND2X0_RVT U6957 ( .A1(n7675), .A2(n7716), .Y(n7715) );
  NAND2X0_RVT U6958 ( .A1(n7717), .A2(n7718), .Y(n7716) );
  NAND2X0_RVT U6959 ( .A1(n7694), .A2(n5022), .Y(n7718) );
  NAND2X0_RVT U6960 ( .A1(n7678), .A2(n5021), .Y(n7717) );
  NAND2X0_RVT U6961 ( .A1(n7679), .A2(n7719), .Y(n7714) );
  NAND2X0_RVT U6962 ( .A1(n7681), .A2(n7720), .Y(n7713) );
  NAND2X0_RVT U6963 ( .A1(n7683), .A2(n7721), .Y(n7712) );
  NAND2X0_RVT U6964 ( .A1(n7722), .A2(n7723), .Y(n7597) );
  NAND2X0_RVT U6965 ( .A1(n7581), .A2(n7579), .Y(n7723) );
  AND2X1_RVT U6966 ( .A1(n7192), .A2(n4984), .Y(n7581) );
  NAND2X0_RVT U6967 ( .A1(n7579), .A2(n7580), .Y(n7722) );
  NAND4X0_RVT U6968 ( .A1(n7724), .A2(n7725), .A3(n7726), .A4(n7727), .Y(n7580) );
  NAND2X0_RVT U6969 ( .A1(n7675), .A2(n7728), .Y(n7727) );
  NAND2X0_RVT U6970 ( .A1(n877), .A2(n7729), .Y(n7728) );
  NAND2X0_RVT U6971 ( .A1(n7678), .A2(n5015), .Y(n7729) );
  NAND2X0_RVT U6972 ( .A1(n7679), .A2(n7730), .Y(n7726) );
  NAND2X0_RVT U6973 ( .A1(n7681), .A2(n7731), .Y(n7725) );
  NAND2X0_RVT U6974 ( .A1(n7683), .A2(n7732), .Y(n7724) );
  NAND2X0_RVT U6975 ( .A1(n7733), .A2(n7734), .Y(n7579) );
  NAND2X0_RVT U6976 ( .A1(n7563), .A2(n7561), .Y(n7734) );
  AND2X1_RVT U6977 ( .A1(n7192), .A2(n4985), .Y(n7563) );
  NAND2X0_RVT U6978 ( .A1(n7561), .A2(n7562), .Y(n7733) );
  NAND4X0_RVT U6979 ( .A1(n7735), .A2(n7736), .A3(n7737), .A4(n7738), .Y(n7562) );
  NAND2X0_RVT U6980 ( .A1(n7675), .A2(n7739), .Y(n7738) );
  NAND2X0_RVT U6981 ( .A1(n7740), .A2(n7741), .Y(n7739) );
  NAND2X0_RVT U6982 ( .A1(n7694), .A2(n5009), .Y(n7741) );
  NAND2X0_RVT U6983 ( .A1(n7678), .A2(n5008), .Y(n7740) );
  NAND2X0_RVT U6984 ( .A1(n7679), .A2(n7742), .Y(n7737) );
  NAND2X0_RVT U6985 ( .A1(n7681), .A2(n7743), .Y(n7736) );
  NAND2X0_RVT U6986 ( .A1(n7683), .A2(n7744), .Y(n7735) );
  AND2X1_RVT U6987 ( .A1(n7745), .A2(n7543), .Y(n7561) );
  NAND4X0_RVT U6988 ( .A1(n7746), .A2(n7747), .A3(n7748), .A4(n7749), .Y(n7543) );
  NAND2X0_RVT U6989 ( .A1(n7683), .A2(n7750), .Y(n7749) );
  AND2X1_RVT U6990 ( .A1(n7751), .A2(n7752), .Y(n7748) );
  NAND2X0_RVT U6991 ( .A1(n7679), .A2(n7753), .Y(n7752) );
  NAND2X0_RVT U6992 ( .A1(n7681), .A2(n7754), .Y(n7751) );
  NAND2X0_RVT U6993 ( .A1(n7675), .A2(n7755), .Y(n7747) );
  NAND2X0_RVT U6994 ( .A1(n7192), .A2(n4990), .Y(n7746) );
  NAND2X0_RVT U6995 ( .A1(n7544), .A2(n7545), .Y(n7745) );
  NAND2X0_RVT U6996 ( .A1(n7527), .A2(n7528), .Y(n7545) );
  NAND4X0_RVT U6997 ( .A1(n7756), .A2(n7757), .A3(n7758), .A4(n7759), .Y(n7528) );
  NAND2X0_RVT U6998 ( .A1(n7683), .A2(n7680), .Y(n7759) );
  AND2X1_RVT U6999 ( .A1(n7760), .A2(n7761), .Y(n7758) );
  NAND2X0_RVT U7000 ( .A1(n7679), .A2(n7762), .Y(n7761) );
  NAND2X0_RVT U7001 ( .A1(n7681), .A2(n7684), .Y(n7760) );
  NAND2X0_RVT U7002 ( .A1(n7675), .A2(n7682), .Y(n7757) );
  NAND3X0_RVT U7003 ( .A1(n7763), .A2(n7764), .A3(n7765), .Y(n7682) );
  NAND2X0_RVT U7004 ( .A1(n7766), .A2(n5111), .Y(n7765) );
  NAND2X0_RVT U7005 ( .A1(n7694), .A2(n5041), .Y(n7764) );
  NAND2X0_RVT U7006 ( .A1(n7678), .A2(n5040), .Y(n7763) );
  NAND2X0_RVT U7007 ( .A1(n7192), .A2(n4991), .Y(n7756) );
  AND3X1_RVT U7008 ( .A1(n7512), .A2(n7496), .A3(n7495), .Y(n7527) );
  AND3X1_RVT U7009 ( .A1(n7480), .A2(n7464), .A3(n7463), .Y(n7495) );
  AND3X1_RVT U7010 ( .A1(n7448), .A2(n7432), .A3(n7431), .Y(n7463) );
  NOR2X0_RVT U7011 ( .A1(n7128), .A2(n9538), .Y(n7431) );
  OR2X1_RVT U7012 ( .A1(n7123), .A2(n9539), .Y(n7128) );
  OR2X1_RVT U7013 ( .A1(n7118), .A2(n9540), .Y(n7123) );
  OR2X1_RVT U7014 ( .A1(n7113), .A2(n9541), .Y(n7118) );
  OR2X1_RVT U7015 ( .A1(n7108), .A2(n9542), .Y(n7113) );
  NAND2X0_RVT U7016 ( .A1(n7102), .A2(n7103), .Y(n7108) );
  AND2X1_RVT U7017 ( .A1(n7192), .A2(n4966), .Y(n7103) );
  NOR2X0_RVT U7018 ( .A1(n7097), .A2(n9515), .Y(n7102) );
  OR2X1_RVT U7019 ( .A1(n7092), .A2(n9516), .Y(n7097) );
  OR2X1_RVT U7020 ( .A1(n7087), .A2(n9517), .Y(n7092) );
  OR2X1_RVT U7021 ( .A1(n7082), .A2(n9518), .Y(n7087) );
  OR2X1_RVT U7022 ( .A1(n7077), .A2(n9519), .Y(n7082) );
  OR2X1_RVT U7023 ( .A1(n7072), .A2(n9520), .Y(n7077) );
  OR2X1_RVT U7024 ( .A1(n7067), .A2(n9522), .Y(n7072) );
  OR2X1_RVT U7025 ( .A1(n7062), .A2(n9533), .Y(n7067) );
  NAND2X0_RVT U7026 ( .A1(n4911), .A2(n4964), .Y(n7062) );
  NAND4X0_RVT U7027 ( .A1(n7767), .A2(n7768), .A3(n7769), .A4(n7770), .Y(n7432) );
  NAND2X0_RVT U7028 ( .A1(n7683), .A2(n7771), .Y(n7770) );
  AND2X1_RVT U7029 ( .A1(n7772), .A2(n7773), .Y(n7769) );
  NAND2X0_RVT U7030 ( .A1(n7679), .A2(n7774), .Y(n7773) );
  NAND2X0_RVT U7031 ( .A1(n7681), .A2(n7775), .Y(n7772) );
  NAND2X0_RVT U7032 ( .A1(n7675), .A2(n7776), .Y(n7768) );
  NAND2X0_RVT U7033 ( .A1(n7192), .A2(n4986), .Y(n7767) );
  NAND4X0_RVT U7034 ( .A1(n7777), .A2(n7778), .A3(n7779), .A4(n7780), .Y(n7448) );
  NAND2X0_RVT U7035 ( .A1(n7683), .A2(n7742), .Y(n7780) );
  AND2X1_RVT U7036 ( .A1(n7781), .A2(n7782), .Y(n7779) );
  NAND2X0_RVT U7037 ( .A1(n7679), .A2(n7783), .Y(n7782) );
  NAND2X0_RVT U7038 ( .A1(n7681), .A2(n7744), .Y(n7781) );
  NAND2X0_RVT U7039 ( .A1(n7675), .A2(n7743), .Y(n7778) );
  NAND3X0_RVT U7040 ( .A1(n7784), .A2(n7785), .A3(n7786), .Y(n7743) );
  NAND2X0_RVT U7041 ( .A1(n7766), .A2(n5112), .Y(n7786) );
  NAND2X0_RVT U7042 ( .A1(n7694), .A2(n5007), .Y(n7785) );
  NAND2X0_RVT U7043 ( .A1(n7678), .A2(n5006), .Y(n7784) );
  NAND2X0_RVT U7044 ( .A1(n7192), .A2(n4987), .Y(n7777) );
  NAND4X0_RVT U7045 ( .A1(n7787), .A2(n7788), .A3(n7789), .A4(n7790), .Y(n7464) );
  NAND2X0_RVT U7046 ( .A1(n7683), .A2(n7730), .Y(n7790) );
  AND2X1_RVT U7047 ( .A1(n7791), .A2(n7792), .Y(n7789) );
  NAND2X0_RVT U7048 ( .A1(n7679), .A2(n7793), .Y(n7792) );
  NAND2X0_RVT U7049 ( .A1(n7681), .A2(n7732), .Y(n7791) );
  NAND2X0_RVT U7050 ( .A1(n7675), .A2(n7731), .Y(n7788) );
  NAND3X0_RVT U7051 ( .A1(n7794), .A2(n7795), .A3(n7796), .Y(n7731) );
  NAND2X0_RVT U7052 ( .A1(n7766), .A2(n5113), .Y(n7796) );
  NAND2X0_RVT U7053 ( .A1(n7694), .A2(n5014), .Y(n7795) );
  NAND2X0_RVT U7054 ( .A1(n7678), .A2(n5013), .Y(n7794) );
  NAND2X0_RVT U7055 ( .A1(n7192), .A2(n4992), .Y(n7787) );
  NAND4X0_RVT U7056 ( .A1(n7797), .A2(n7798), .A3(n7799), .A4(n7800), .Y(n7480) );
  NAND2X0_RVT U7057 ( .A1(n7683), .A2(n7719), .Y(n7800) );
  AND2X1_RVT U7058 ( .A1(n7801), .A2(n7802), .Y(n7799) );
  NAND2X0_RVT U7059 ( .A1(n7679), .A2(n7803), .Y(n7802) );
  NAND2X0_RVT U7060 ( .A1(n7681), .A2(n7721), .Y(n7801) );
  NAND2X0_RVT U7061 ( .A1(n7675), .A2(n7720), .Y(n7798) );
  NAND3X0_RVT U7062 ( .A1(n7804), .A2(n7805), .A3(n7806), .Y(n7720) );
  NAND2X0_RVT U7063 ( .A1(n7766), .A2(n5114), .Y(n7806) );
  NAND2X0_RVT U7064 ( .A1(n7694), .A2(n5020), .Y(n7805) );
  NAND2X0_RVT U7065 ( .A1(n7678), .A2(n5019), .Y(n7804) );
  NAND2X0_RVT U7066 ( .A1(n7192), .A2(n4993), .Y(n7797) );
  NAND4X0_RVT U7067 ( .A1(n7807), .A2(n7808), .A3(n7809), .A4(n7810), .Y(n7496) );
  NAND2X0_RVT U7068 ( .A1(n7683), .A2(n7707), .Y(n7810) );
  AND2X1_RVT U7069 ( .A1(n7811), .A2(n7812), .Y(n7809) );
  NAND2X0_RVT U7070 ( .A1(n7679), .A2(n7813), .Y(n7812) );
  NAND2X0_RVT U7071 ( .A1(n7681), .A2(n7709), .Y(n7811) );
  NAND2X0_RVT U7072 ( .A1(n7675), .A2(n7708), .Y(n7808) );
  NAND3X0_RVT U7073 ( .A1(n7814), .A2(n7815), .A3(n7816), .Y(n7708) );
  NAND2X0_RVT U7074 ( .A1(n7766), .A2(n5115), .Y(n7816) );
  NAND2X0_RVT U7075 ( .A1(n7694), .A2(n5027), .Y(n7815) );
  NAND2X0_RVT U7076 ( .A1(n7678), .A2(n5026), .Y(n7814) );
  NAND2X0_RVT U7077 ( .A1(n7192), .A2(n4994), .Y(n7807) );
  NAND4X0_RVT U7078 ( .A1(n7817), .A2(n7818), .A3(n7819), .A4(n7820), .Y(n7512) );
  NAND2X0_RVT U7079 ( .A1(n7683), .A2(n7695), .Y(n7820) );
  AND2X1_RVT U7080 ( .A1(n7821), .A2(n7822), .Y(n7819) );
  NAND2X0_RVT U7081 ( .A1(n7679), .A2(n7823), .Y(n7822) );
  NAND2X0_RVT U7082 ( .A1(n7681), .A2(n7697), .Y(n7821) );
  NAND2X0_RVT U7083 ( .A1(n7675), .A2(n7696), .Y(n7818) );
  NAND3X0_RVT U7084 ( .A1(n7824), .A2(n7825), .A3(n7826), .Y(n7696) );
  NAND2X0_RVT U7085 ( .A1(n7766), .A2(n5116), .Y(n7826) );
  NAND2X0_RVT U7086 ( .A1(n7694), .A2(n5034), .Y(n7825) );
  NAND2X0_RVT U7087 ( .A1(n7678), .A2(n5033), .Y(n7824) );
  NAND2X0_RVT U7088 ( .A1(n7192), .A2(n4995), .Y(n7817) );
  AND4X1_RVT U7089 ( .A1(n7827), .A2(n7828), .A3(n7829), .A4(n7830), .Y(n7544)
         );
  NAND2X0_RVT U7090 ( .A1(n7675), .A2(n7831), .Y(n7830) );
  NAND2X0_RVT U7091 ( .A1(n7832), .A2(n7833), .Y(n7831) );
  NAND2X0_RVT U7092 ( .A1(n7694), .A2(n5002), .Y(n7833) );
  NAND2X0_RVT U7093 ( .A1(n7678), .A2(n5001), .Y(n7832) );
  NAND2X0_RVT U7094 ( .A1(n7679), .A2(n7771), .Y(n7829) );
  NAND2X0_RVT U7095 ( .A1(n7681), .A2(n7776), .Y(n7828) );
  NAND3X0_RVT U7096 ( .A1(n7834), .A2(n7835), .A3(n7836), .Y(n7776) );
  NAND2X0_RVT U7097 ( .A1(n7766), .A2(n5117), .Y(n7836) );
  NAND2X0_RVT U7098 ( .A1(n7694), .A2(n5000), .Y(n7835) );
  NAND2X0_RVT U7099 ( .A1(n7678), .A2(n4999), .Y(n7834) );
  NAND2X0_RVT U7100 ( .A1(n7683), .A2(n7775), .Y(n7827) );
  NAND4X0_RVT U7101 ( .A1(n7837), .A2(n7838), .A3(n7839), .A4(n7840), .Y(n7668) );
  NAND2X0_RVT U7102 ( .A1(n7679), .A2(n7750), .Y(n7840) );
  AND2X1_RVT U7103 ( .A1(n7841), .A2(n7842), .Y(n7679) );
  AND2X1_RVT U7104 ( .A1(n7843), .A2(n7196), .Y(n7839) );
  NAND2X0_RVT U7105 ( .A1(n7192), .A2(n4988), .Y(n7196) );
  NAND2X0_RVT U7106 ( .A1(n7675), .A2(n7845), .Y(n7843) );
  NAND2X0_RVT U7107 ( .A1(n7846), .A2(n7847), .Y(n7845) );
  NAND2X0_RVT U7108 ( .A1(n7694), .A2(n5050), .Y(n7847) );
  NAND2X0_RVT U7109 ( .A1(n7678), .A2(n5051), .Y(n7846) );
  AND2X1_RVT U7110 ( .A1(n7841), .A2(n7848), .Y(n7675) );
  NAND2X0_RVT U7111 ( .A1(n7681), .A2(n7755), .Y(n7838) );
  NAND3X0_RVT U7112 ( .A1(n7849), .A2(n7850), .A3(n7851), .Y(n7755) );
  NAND2X0_RVT U7113 ( .A1(n7766), .A2(n5048), .Y(n7851) );
  NAND2X0_RVT U7114 ( .A1(n7694), .A2(n5046), .Y(n7850) );
  NAND2X0_RVT U7115 ( .A1(n7678), .A2(n5047), .Y(n7849) );
  AND2X1_RVT U7116 ( .A1(n7841), .A2(n7852), .Y(n7681) );
  NAND2X0_RVT U7117 ( .A1(n7683), .A2(n7754), .Y(n7837) );
  AND2X1_RVT U7118 ( .A1(n7841), .A2(n7853), .Y(n7683) );
  INVX0_RVT U7119 ( .A(n6497), .Y(n7841) );
  NAND2X0_RVT U7120 ( .A1(n7218), .A2(rEIP[30]), .Y(n7654) );
  NAND4X0_RVT U7121 ( .A1(n7854), .A2(n7855), .A3(n7856), .A4(n7857), .Y(n4589) );
  AND3X1_RVT U7122 ( .A1(n7858), .A2(n7859), .A3(n7860), .Y(n7857) );
  NAND2X0_RVT U7123 ( .A1(n7215), .A2(n5086), .Y(n7860) );
  NAND2X0_RVT U7124 ( .A1(n7861), .A2(n7214), .Y(n7859) );
  NAND2X0_RVT U7125 ( .A1(n7864), .A2(n7865), .Y(n7862) );
  NAND2X0_RVT U7126 ( .A1(n7218), .A2(rEIP[31]), .Y(n7858) );
  NAND2X0_RVT U7127 ( .A1(n7212), .A2(n4958), .Y(n7856) );
  NAND2X0_RVT U7128 ( .A1(n7867), .A2(n7868), .Y(n7866) );
  NAND3X0_RVT U7129 ( .A1(n7046), .A2(n7869), .A3(n7864), .Y(n7868) );
  NAND2X0_RVT U7130 ( .A1(n5272), .A2(n7870), .Y(n7867) );
  NAND2X0_RVT U7131 ( .A1(n7871), .A2(n5271), .Y(n7870) );
  NAND2X0_RVT U7132 ( .A1(n7667), .A2(n7666), .Y(n7855) );
  AND2X1_RVT U7133 ( .A1(n7649), .A2(n7648), .Y(n7666) );
  AND2X1_RVT U7134 ( .A1(n7631), .A2(n7630), .Y(n7648) );
  AND2X1_RVT U7135 ( .A1(n7613), .A2(n7612), .Y(n7630) );
  AND2X1_RVT U7136 ( .A1(n7595), .A2(n7594), .Y(n7612) );
  AND2X1_RVT U7137 ( .A1(n7577), .A2(n7576), .Y(n7594) );
  AND2X1_RVT U7138 ( .A1(n7559), .A2(n7558), .Y(n7576) );
  AND2X1_RVT U7139 ( .A1(n7542), .A2(n7541), .Y(n7558) );
  AND2X1_RVT U7140 ( .A1(n7526), .A2(n7525), .Y(n7541) );
  AND2X1_RVT U7141 ( .A1(n7510), .A2(n7509), .Y(n7525) );
  AND2X1_RVT U7142 ( .A1(n7494), .A2(n7493), .Y(n7509) );
  AND2X1_RVT U7143 ( .A1(n7478), .A2(n7477), .Y(n7493) );
  AND2X1_RVT U7144 ( .A1(n7462), .A2(n7461), .Y(n7477) );
  AND2X1_RVT U7145 ( .A1(n7446), .A2(n7445), .Y(n7461) );
  AND2X1_RVT U7146 ( .A1(n7429), .A2(n7428), .Y(n7445) );
  NOR2X0_RVT U7147 ( .A1(n7415), .A2(n7414), .Y(n7428) );
  OR2X1_RVT U7148 ( .A1(n7404), .A2(n7403), .Y(n7414) );
  OR2X1_RVT U7149 ( .A1(n7393), .A2(n7392), .Y(n7403) );
  OR2X1_RVT U7150 ( .A1(n7382), .A2(n7381), .Y(n7392) );
  OR2X1_RVT U7151 ( .A1(n7371), .A2(n7370), .Y(n7381) );
  OR2X1_RVT U7152 ( .A1(n7360), .A2(n7359), .Y(n7370) );
  OR2X1_RVT U7153 ( .A1(n7349), .A2(n7348), .Y(n7359) );
  OR2X1_RVT U7154 ( .A1(n7338), .A2(n7337), .Y(n7348) );
  OR2X1_RVT U7155 ( .A1(n7327), .A2(n7326), .Y(n7337) );
  OR2X1_RVT U7156 ( .A1(n7316), .A2(n7315), .Y(n7326) );
  OR2X1_RVT U7157 ( .A1(n7305), .A2(n7304), .Y(n7315) );
  NAND2X0_RVT U7158 ( .A1(n7293), .A2(n7294), .Y(n7304) );
  AND2X1_RVT U7159 ( .A1(n7282), .A2(n7283), .Y(n7294) );
  AND2X1_RVT U7160 ( .A1(n7249), .A2(n7250), .Y(n7283) );
  AND2X1_RVT U7161 ( .A1(n7234), .A2(n7233), .Y(n7250) );
  XNOR2X1_RVT U7162 ( .A1(n7872), .A2(n7217), .Y(n7233) );
  NAND2X0_RVT U7163 ( .A1(n7442), .A2(n7873), .Y(n7872) );
  NAND2X0_RVT U7164 ( .A1(n7232), .A2(n7874), .Y(n7873) );
  NAND2X0_RVT U7165 ( .A1(n7875), .A2(Datai[1]), .Y(n7442) );
  AND2X1_RVT U7166 ( .A1(n7216), .A2(n7876), .Y(n7234) );
  XNOR2X1_RVT U7167 ( .A1(n7877), .A2(n7217), .Y(n7216) );
  NAND2X0_RVT U7168 ( .A1(n7425), .A2(n7878), .Y(n7877) );
  NAND2X0_RVT U7169 ( .A1(n7213), .A2(n7874), .Y(n7878) );
  NAND2X0_RVT U7170 ( .A1(n7875), .A2(Datai[0]), .Y(n7425) );
  XNOR2X1_RVT U7171 ( .A1(n7879), .A2(n7217), .Y(n7249) );
  NAND2X0_RVT U7172 ( .A1(n7458), .A2(n7880), .Y(n7879) );
  NAND2X0_RVT U7173 ( .A1(n7248), .A2(n7874), .Y(n7880) );
  NAND2X0_RVT U7174 ( .A1(n7875), .A2(Datai[2]), .Y(n7458) );
  XNOR2X1_RVT U7175 ( .A1(n7881), .A2(n7217), .Y(n7282) );
  NAND2X0_RVT U7176 ( .A1(n7474), .A2(n7882), .Y(n7881) );
  NAND2X0_RVT U7177 ( .A1(n7281), .A2(n7874), .Y(n7882) );
  NAND2X0_RVT U7178 ( .A1(n7875), .A2(Datai[3]), .Y(n7474) );
  XNOR2X1_RVT U7179 ( .A1(n7883), .A2(n7217), .Y(n7293) );
  NAND2X0_RVT U7180 ( .A1(n7490), .A2(n7884), .Y(n7883) );
  NAND2X0_RVT U7181 ( .A1(n7292), .A2(n7874), .Y(n7884) );
  NAND2X0_RVT U7182 ( .A1(n7875), .A2(Datai[4]), .Y(n7490) );
  XOR2X1_RVT U7183 ( .A1(n7885), .A2(n7217), .Y(n7305) );
  NAND2X0_RVT U7184 ( .A1(n7506), .A2(n7886), .Y(n7885) );
  NAND2X0_RVT U7185 ( .A1(n7303), .A2(n7874), .Y(n7886) );
  NAND2X0_RVT U7186 ( .A1(n7875), .A2(Datai[5]), .Y(n7506) );
  XOR2X1_RVT U7187 ( .A1(n7887), .A2(n7217), .Y(n7316) );
  NAND2X0_RVT U7188 ( .A1(n7522), .A2(n7888), .Y(n7887) );
  NAND2X0_RVT U7189 ( .A1(n7314), .A2(n7874), .Y(n7888) );
  NAND2X0_RVT U7190 ( .A1(n7875), .A2(Datai[6]), .Y(n7522) );
  XOR2X1_RVT U7191 ( .A1(n7889), .A2(n7217), .Y(n7327) );
  NAND2X0_RVT U7192 ( .A1(n7538), .A2(n7890), .Y(n7889) );
  NAND2X0_RVT U7193 ( .A1(n7325), .A2(n7874), .Y(n7890) );
  NAND2X0_RVT U7194 ( .A1(n7875), .A2(Datai[7]), .Y(n7538) );
  XOR2X1_RVT U7195 ( .A1(n7891), .A2(n7217), .Y(n7338) );
  NAND2X0_RVT U7196 ( .A1(n7555), .A2(n7892), .Y(n7891) );
  NAND2X0_RVT U7197 ( .A1(n7336), .A2(n7874), .Y(n7892) );
  NAND2X0_RVT U7198 ( .A1(Datai[8]), .A2(n7875), .Y(n7555) );
  XOR2X1_RVT U7199 ( .A1(n7893), .A2(n7217), .Y(n7349) );
  NAND2X0_RVT U7200 ( .A1(n7573), .A2(n7894), .Y(n7893) );
  NAND2X0_RVT U7201 ( .A1(n7347), .A2(n7874), .Y(n7894) );
  NAND2X0_RVT U7202 ( .A1(Datai[9]), .A2(n7875), .Y(n7573) );
  XOR2X1_RVT U7203 ( .A1(n7895), .A2(n7217), .Y(n7360) );
  NAND2X0_RVT U7204 ( .A1(n7591), .A2(n7896), .Y(n7895) );
  NAND2X0_RVT U7205 ( .A1(n7358), .A2(n7874), .Y(n7896) );
  NAND2X0_RVT U7206 ( .A1(Datai[10]), .A2(n7875), .Y(n7591) );
  XOR2X1_RVT U7207 ( .A1(n7897), .A2(n7217), .Y(n7371) );
  NAND2X0_RVT U7208 ( .A1(n7609), .A2(n7898), .Y(n7897) );
  NAND2X0_RVT U7209 ( .A1(n7369), .A2(n7874), .Y(n7898) );
  NAND2X0_RVT U7210 ( .A1(Datai[11]), .A2(n7875), .Y(n7609) );
  XOR2X1_RVT U7211 ( .A1(n7899), .A2(n7217), .Y(n7382) );
  NAND2X0_RVT U7212 ( .A1(n7627), .A2(n7900), .Y(n7899) );
  NAND2X0_RVT U7213 ( .A1(n7380), .A2(n7874), .Y(n7900) );
  NAND2X0_RVT U7214 ( .A1(Datai[12]), .A2(n7875), .Y(n7627) );
  XOR2X1_RVT U7215 ( .A1(n7901), .A2(n7217), .Y(n7393) );
  NAND2X0_RVT U7216 ( .A1(n7645), .A2(n7902), .Y(n7901) );
  NAND2X0_RVT U7217 ( .A1(n7391), .A2(n7874), .Y(n7902) );
  NAND2X0_RVT U7218 ( .A1(Datai[13]), .A2(n7875), .Y(n7645) );
  XOR2X1_RVT U7219 ( .A1(n7903), .A2(n7217), .Y(n7404) );
  NAND2X0_RVT U7220 ( .A1(n7663), .A2(n7904), .Y(n7903) );
  NAND2X0_RVT U7221 ( .A1(n7402), .A2(n7874), .Y(n7904) );
  NAND2X0_RVT U7222 ( .A1(Datai[14]), .A2(n7875), .Y(n7663) );
  XOR2X1_RVT U7223 ( .A1(n7905), .A2(n7217), .Y(n7415) );
  NAND2X0_RVT U7224 ( .A1(n7906), .A2(n7907), .Y(n7905) );
  NAND2X0_RVT U7225 ( .A1(n7413), .A2(n7874), .Y(n7907) );
  OR2X1_RVT U7226 ( .A1(n7430), .A2(n7876), .Y(n7874) );
  INVX0_RVT U7227 ( .A(n7217), .Y(n7876) );
  NAND2X0_RVT U7228 ( .A1(Datai[15]), .A2(n7875), .Y(n7906) );
  NOR2X0_RVT U7229 ( .A1(n7217), .A2(n7424), .Y(n7429) );
  NOR2X0_RVT U7230 ( .A1(n7217), .A2(n7441), .Y(n7446) );
  NOR2X0_RVT U7231 ( .A1(n7217), .A2(n7457), .Y(n7462) );
  NOR2X0_RVT U7232 ( .A1(n7217), .A2(n7473), .Y(n7478) );
  NOR2X0_RVT U7233 ( .A1(n7217), .A2(n7488), .Y(n7494) );
  NOR2X0_RVT U7234 ( .A1(n7217), .A2(n7504), .Y(n7510) );
  NOR2X0_RVT U7235 ( .A1(n7217), .A2(n7520), .Y(n7526) );
  NOR2X0_RVT U7236 ( .A1(n7217), .A2(n7536), .Y(n7542) );
  NOR2X0_RVT U7237 ( .A1(n7217), .A2(n7553), .Y(n7559) );
  NOR2X0_RVT U7238 ( .A1(n7217), .A2(n7571), .Y(n7577) );
  NOR2X0_RVT U7239 ( .A1(n7217), .A2(n7589), .Y(n7595) );
  NOR2X0_RVT U7240 ( .A1(n7217), .A2(n7607), .Y(n7613) );
  NOR2X0_RVT U7241 ( .A1(n7217), .A2(n7625), .Y(n7631) );
  NOR2X0_RVT U7242 ( .A1(n7217), .A2(n7643), .Y(n7649) );
  NOR2X0_RVT U7243 ( .A1(n7217), .A2(n7661), .Y(n7667) );
  NAND3X0_RVT U7244 ( .A1(n7909), .A2(n7210), .A3(n7910), .Y(n7854) );
  INVX0_RVT U7245 ( .A(n7863), .Y(n7207) );
  NAND2X0_RVT U7246 ( .A1(n5265), .A2(n7865), .Y(n7863) );
  NAND2X0_RVT U7247 ( .A1(n7009), .A2(n7911), .Y(n6755) );
  NAND2X0_RVT U7248 ( .A1(n7912), .A2(n6756), .Y(n7911) );
  NAND3X0_RVT U7249 ( .A1(n4925), .A2(n4969), .A3(n6760), .Y(n6446) );
  NAND2X0_RVT U7250 ( .A1(n7913), .A2(n7914), .Y(n4588) );
  XNOR2X1_RVT U7251 ( .A1(n7915), .A2(n7916), .Y(n7914) );
  NAND2X0_RVT U7252 ( .A1(n5276), .A2(Address[0]), .Y(n7913) );
  NAND2X0_RVT U7253 ( .A1(n7917), .A2(n7918), .Y(n4587) );
  XOR2X1_RVT U7254 ( .A1(n7919), .A2(n7920), .Y(n7918) );
  NAND2X0_RVT U7255 ( .A1(n7915), .A2(n7916), .Y(n7920) );
  NAND2X0_RVT U7256 ( .A1(n5276), .A2(Address[1]), .Y(n7917) );
  NAND2X0_RVT U7257 ( .A1(n7921), .A2(n7922), .Y(n4586) );
  XNOR2X1_RVT U7258 ( .A1(n7923), .A2(n7924), .Y(n7922) );
  NAND2X0_RVT U7259 ( .A1(n5276), .A2(Address[2]), .Y(n7921) );
  NAND2X0_RVT U7260 ( .A1(n7925), .A2(n7926), .Y(n4585) );
  XOR2X1_RVT U7261 ( .A1(n7927), .A2(n7928), .Y(n7926) );
  NAND2X0_RVT U7262 ( .A1(n7923), .A2(n7924), .Y(n7928) );
  NAND2X0_RVT U7263 ( .A1(n5276), .A2(Address[3]), .Y(n7925) );
  NAND2X0_RVT U7264 ( .A1(n7929), .A2(n7930), .Y(n4584) );
  XNOR2X1_RVT U7265 ( .A1(n7931), .A2(n7932), .Y(n7930) );
  NAND2X0_RVT U7266 ( .A1(n5276), .A2(Address[4]), .Y(n7929) );
  NAND2X0_RVT U7267 ( .A1(n7933), .A2(n7934), .Y(n4583) );
  XOR2X1_RVT U7268 ( .A1(n7935), .A2(n7936), .Y(n7934) );
  NAND2X0_RVT U7269 ( .A1(n7931), .A2(n7932), .Y(n7936) );
  NAND2X0_RVT U7270 ( .A1(n5276), .A2(Address[5]), .Y(n7933) );
  NAND2X0_RVT U7271 ( .A1(n7937), .A2(n7938), .Y(n4582) );
  XNOR2X1_RVT U7272 ( .A1(n7939), .A2(n7940), .Y(n7938) );
  NAND2X0_RVT U7273 ( .A1(n5276), .A2(Address[6]), .Y(n7937) );
  NAND2X0_RVT U7274 ( .A1(n7941), .A2(n7942), .Y(n4581) );
  XOR2X1_RVT U7275 ( .A1(n7943), .A2(n7944), .Y(n7942) );
  NAND2X0_RVT U7276 ( .A1(n7939), .A2(n7940), .Y(n7944) );
  NAND2X0_RVT U7277 ( .A1(n5276), .A2(Address[7]), .Y(n7941) );
  NAND2X0_RVT U7278 ( .A1(n7945), .A2(n7946), .Y(n4580) );
  XNOR2X1_RVT U7279 ( .A1(n7947), .A2(n7948), .Y(n7946) );
  NAND2X0_RVT U7280 ( .A1(n5276), .A2(Address[8]), .Y(n7945) );
  NAND2X0_RVT U7281 ( .A1(n7949), .A2(n7950), .Y(n4579) );
  XOR2X1_RVT U7282 ( .A1(n7951), .A2(n7952), .Y(n7950) );
  NAND2X0_RVT U7283 ( .A1(n7947), .A2(n7948), .Y(n7952) );
  NAND2X0_RVT U7284 ( .A1(n5276), .A2(Address[9]), .Y(n7949) );
  NAND2X0_RVT U7285 ( .A1(n7953), .A2(n7954), .Y(n4578) );
  XNOR2X1_RVT U7286 ( .A1(n7955), .A2(n7956), .Y(n7954) );
  NAND2X0_RVT U7287 ( .A1(n5276), .A2(Address[10]), .Y(n7953) );
  NAND2X0_RVT U7288 ( .A1(n7957), .A2(n7958), .Y(n4577) );
  XOR2X1_RVT U7289 ( .A1(n7959), .A2(n7960), .Y(n7958) );
  NAND2X0_RVT U7290 ( .A1(n7955), .A2(n7956), .Y(n7960) );
  NAND2X0_RVT U7291 ( .A1(n5276), .A2(Address[11]), .Y(n7957) );
  NAND2X0_RVT U7292 ( .A1(n7961), .A2(n7962), .Y(n4576) );
  XNOR2X1_RVT U7293 ( .A1(n7963), .A2(n7964), .Y(n7962) );
  NAND2X0_RVT U7294 ( .A1(n5276), .A2(Address[12]), .Y(n7961) );
  NAND2X0_RVT U7295 ( .A1(n7965), .A2(n7966), .Y(n4575) );
  XOR2X1_RVT U7296 ( .A1(n7967), .A2(n7968), .Y(n7966) );
  NAND2X0_RVT U7297 ( .A1(n7963), .A2(n7964), .Y(n7968) );
  NAND2X0_RVT U7298 ( .A1(n5276), .A2(Address[13]), .Y(n7965) );
  NAND2X0_RVT U7299 ( .A1(n7969), .A2(n7970), .Y(n4574) );
  XNOR2X1_RVT U7300 ( .A1(n7971), .A2(n7972), .Y(n7970) );
  NAND2X0_RVT U7301 ( .A1(n5276), .A2(Address[14]), .Y(n7969) );
  NAND2X0_RVT U7302 ( .A1(n7973), .A2(n7974), .Y(n4573) );
  XOR2X1_RVT U7303 ( .A1(n7975), .A2(n7976), .Y(n7974) );
  NAND2X0_RVT U7304 ( .A1(n7971), .A2(n7972), .Y(n7976) );
  NAND2X0_RVT U7305 ( .A1(n5276), .A2(Address[15]), .Y(n7973) );
  NAND2X0_RVT U7306 ( .A1(n7977), .A2(n7978), .Y(n4572) );
  XNOR2X1_RVT U7307 ( .A1(n7979), .A2(n7980), .Y(n7978) );
  NAND2X0_RVT U7308 ( .A1(n5276), .A2(Address[16]), .Y(n7977) );
  NAND2X0_RVT U7309 ( .A1(n7981), .A2(n7982), .Y(n4571) );
  XOR2X1_RVT U7310 ( .A1(n7983), .A2(n7984), .Y(n7982) );
  NAND2X0_RVT U7311 ( .A1(n7979), .A2(n7980), .Y(n7984) );
  NAND2X0_RVT U7312 ( .A1(n5276), .A2(Address[17]), .Y(n7981) );
  NAND2X0_RVT U7313 ( .A1(n7985), .A2(n7986), .Y(n4570) );
  XNOR2X1_RVT U7314 ( .A1(n7987), .A2(n7988), .Y(n7986) );
  NAND2X0_RVT U7315 ( .A1(n5276), .A2(Address[18]), .Y(n7985) );
  NAND2X0_RVT U7316 ( .A1(n7989), .A2(n7990), .Y(n4569) );
  XOR2X1_RVT U7317 ( .A1(n7991), .A2(n7992), .Y(n7990) );
  NAND2X0_RVT U7318 ( .A1(n7987), .A2(n7988), .Y(n7992) );
  NAND2X0_RVT U7319 ( .A1(n5276), .A2(Address[19]), .Y(n7989) );
  NAND2X0_RVT U7320 ( .A1(n7993), .A2(n7994), .Y(n4568) );
  XNOR2X1_RVT U7321 ( .A1(n7995), .A2(n7996), .Y(n7994) );
  NAND2X0_RVT U7322 ( .A1(n5276), .A2(Address[20]), .Y(n7993) );
  NAND2X0_RVT U7323 ( .A1(n7997), .A2(n7998), .Y(n4567) );
  XOR2X1_RVT U7324 ( .A1(n7999), .A2(n8000), .Y(n7998) );
  NAND2X0_RVT U7325 ( .A1(n7995), .A2(n7996), .Y(n8000) );
  NAND2X0_RVT U7326 ( .A1(n5276), .A2(Address[21]), .Y(n7997) );
  NAND2X0_RVT U7327 ( .A1(n8001), .A2(n8002), .Y(n4566) );
  XNOR2X1_RVT U7328 ( .A1(n8003), .A2(n8004), .Y(n8002) );
  NAND2X0_RVT U7329 ( .A1(n5276), .A2(Address[22]), .Y(n8001) );
  NAND2X0_RVT U7330 ( .A1(n8005), .A2(n8006), .Y(n4565) );
  XOR2X1_RVT U7331 ( .A1(n8007), .A2(n8008), .Y(n8006) );
  NAND2X0_RVT U7332 ( .A1(n8003), .A2(n8004), .Y(n8008) );
  NAND2X0_RVT U7333 ( .A1(n5276), .A2(Address[23]), .Y(n8005) );
  NAND2X0_RVT U7334 ( .A1(n8009), .A2(n8010), .Y(n4564) );
  XNOR2X1_RVT U7335 ( .A1(n8011), .A2(n8012), .Y(n8010) );
  NAND2X0_RVT U7336 ( .A1(n5276), .A2(Address[24]), .Y(n8009) );
  NAND2X0_RVT U7337 ( .A1(n8013), .A2(n8014), .Y(n4563) );
  XOR2X1_RVT U7338 ( .A1(n8015), .A2(n8016), .Y(n8014) );
  NAND2X0_RVT U7339 ( .A1(n8011), .A2(n8012), .Y(n8016) );
  NAND2X0_RVT U7340 ( .A1(n5276), .A2(Address[25]), .Y(n8013) );
  NAND2X0_RVT U7341 ( .A1(n8017), .A2(n8018), .Y(n4562) );
  XNOR2X1_RVT U7342 ( .A1(n8019), .A2(n8020), .Y(n8018) );
  NAND2X0_RVT U7343 ( .A1(n5276), .A2(Address[26]), .Y(n8017) );
  NAND2X0_RVT U7344 ( .A1(n8021), .A2(n8022), .Y(n4561) );
  XOR2X1_RVT U7345 ( .A1(n8023), .A2(n8024), .Y(n8022) );
  NAND2X0_RVT U7346 ( .A1(n8019), .A2(n8020), .Y(n8024) );
  NAND2X0_RVT U7347 ( .A1(n5276), .A2(Address[27]), .Y(n8021) );
  NAND2X0_RVT U7348 ( .A1(n8025), .A2(n8026), .Y(n4560) );
  XNOR2X1_RVT U7349 ( .A1(n8027), .A2(n8028), .Y(n8026) );
  NAND2X0_RVT U7350 ( .A1(n5276), .A2(Address[28]), .Y(n8025) );
  NAND2X0_RVT U7351 ( .A1(n8029), .A2(n8030), .Y(n4559) );
  XOR2X1_RVT U7352 ( .A1(n8031), .A2(n8032), .Y(n8030) );
  NAND2X0_RVT U7353 ( .A1(n8027), .A2(n8028), .Y(n8032) );
  NAND2X0_RVT U7354 ( .A1(n8033), .A2(n8034), .Y(n8028) );
  NAND2X0_RVT U7355 ( .A1(n8035), .A2(rEIP[29]), .Y(n8034) );
  NAND2X0_RVT U7356 ( .A1(n8036), .A2(rEIP[30]), .Y(n8033) );
  AND3X1_RVT U7357 ( .A1(n8023), .A2(n8020), .A3(n8019), .Y(n8027) );
  AND3X1_RVT U7358 ( .A1(n8015), .A2(n8012), .A3(n8011), .Y(n8019) );
  AND3X1_RVT U7359 ( .A1(n8007), .A2(n8004), .A3(n8003), .Y(n8011) );
  AND3X1_RVT U7360 ( .A1(n7999), .A2(n7996), .A3(n7995), .Y(n8003) );
  AND3X1_RVT U7361 ( .A1(n7991), .A2(n7988), .A3(n7987), .Y(n7995) );
  AND3X1_RVT U7362 ( .A1(n7983), .A2(n7980), .A3(n7979), .Y(n7987) );
  AND3X1_RVT U7363 ( .A1(n7975), .A2(n7972), .A3(n7971), .Y(n7979) );
  AND3X1_RVT U7364 ( .A1(n7967), .A2(n7964), .A3(n7963), .Y(n7971) );
  AND3X1_RVT U7365 ( .A1(n7959), .A2(n7956), .A3(n7955), .Y(n7963) );
  AND3X1_RVT U7366 ( .A1(n7951), .A2(n7948), .A3(n7947), .Y(n7955) );
  AND3X1_RVT U7367 ( .A1(n7943), .A2(n7940), .A3(n7939), .Y(n7947) );
  AND3X1_RVT U7368 ( .A1(n7935), .A2(n7932), .A3(n7931), .Y(n7939) );
  AND3X1_RVT U7369 ( .A1(n7927), .A2(n7924), .A3(n7923), .Y(n7931) );
  AND3X1_RVT U7370 ( .A1(n7919), .A2(n7916), .A3(n7915), .Y(n7923) );
  AND2X1_RVT U7371 ( .A1(rEIP[31]), .A2(n8037), .Y(n7915) );
  NAND2X0_RVT U7372 ( .A1(n8038), .A2(n8039), .Y(n8037) );
  NAND2X0_RVT U7373 ( .A1(rEIP[0]), .A2(n6751), .Y(n8039) );
  NAND2X0_RVT U7374 ( .A1(n8036), .A2(rEIP[1]), .Y(n8038) );
  NAND2X0_RVT U7375 ( .A1(n8040), .A2(n8041), .Y(n7916) );
  NAND2X0_RVT U7376 ( .A1(n8035), .A2(rEIP[1]), .Y(n8041) );
  NAND2X0_RVT U7377 ( .A1(n8036), .A2(rEIP[2]), .Y(n8040) );
  NAND2X0_RVT U7378 ( .A1(n8042), .A2(n8043), .Y(n7919) );
  NAND2X0_RVT U7379 ( .A1(n8035), .A2(rEIP[2]), .Y(n8043) );
  NAND2X0_RVT U7380 ( .A1(n8036), .A2(rEIP[3]), .Y(n8042) );
  NAND2X0_RVT U7381 ( .A1(n8044), .A2(n8045), .Y(n7924) );
  NAND2X0_RVT U7382 ( .A1(n8035), .A2(rEIP[3]), .Y(n8045) );
  NAND2X0_RVT U7383 ( .A1(n8036), .A2(rEIP[4]), .Y(n8044) );
  NAND2X0_RVT U7384 ( .A1(n8046), .A2(n8047), .Y(n7927) );
  NAND2X0_RVT U7385 ( .A1(n8035), .A2(rEIP[4]), .Y(n8047) );
  NAND2X0_RVT U7386 ( .A1(n8036), .A2(rEIP[5]), .Y(n8046) );
  NAND2X0_RVT U7387 ( .A1(n8048), .A2(n8049), .Y(n7932) );
  NAND2X0_RVT U7388 ( .A1(n8035), .A2(rEIP[5]), .Y(n8049) );
  NAND2X0_RVT U7389 ( .A1(n8036), .A2(rEIP[6]), .Y(n8048) );
  NAND2X0_RVT U7390 ( .A1(n8050), .A2(n8051), .Y(n7935) );
  NAND2X0_RVT U7391 ( .A1(n8035), .A2(rEIP[6]), .Y(n8051) );
  NAND2X0_RVT U7392 ( .A1(n8036), .A2(rEIP[7]), .Y(n8050) );
  NAND2X0_RVT U7393 ( .A1(n8052), .A2(n8053), .Y(n7940) );
  NAND2X0_RVT U7394 ( .A1(n8035), .A2(rEIP[7]), .Y(n8053) );
  NAND2X0_RVT U7395 ( .A1(n8036), .A2(rEIP[8]), .Y(n8052) );
  NAND2X0_RVT U7396 ( .A1(n8054), .A2(n8055), .Y(n7943) );
  NAND2X0_RVT U7397 ( .A1(n8035), .A2(rEIP[8]), .Y(n8055) );
  NAND2X0_RVT U7398 ( .A1(n8036), .A2(rEIP[9]), .Y(n8054) );
  NAND2X0_RVT U7399 ( .A1(n8056), .A2(n8057), .Y(n7948) );
  NAND2X0_RVT U7400 ( .A1(n8035), .A2(rEIP[9]), .Y(n8057) );
  NAND2X0_RVT U7401 ( .A1(n8036), .A2(rEIP[10]), .Y(n8056) );
  NAND2X0_RVT U7402 ( .A1(n8058), .A2(n8059), .Y(n7951) );
  NAND2X0_RVT U7403 ( .A1(n8035), .A2(rEIP[10]), .Y(n8059) );
  NAND2X0_RVT U7404 ( .A1(n8036), .A2(rEIP[11]), .Y(n8058) );
  NAND2X0_RVT U7405 ( .A1(n8060), .A2(n8061), .Y(n7956) );
  NAND2X0_RVT U7406 ( .A1(n8035), .A2(rEIP[11]), .Y(n8061) );
  NAND2X0_RVT U7407 ( .A1(n8036), .A2(rEIP[12]), .Y(n8060) );
  NAND2X0_RVT U7408 ( .A1(n8062), .A2(n8063), .Y(n7959) );
  NAND2X0_RVT U7409 ( .A1(n8035), .A2(rEIP[12]), .Y(n8063) );
  NAND2X0_RVT U7410 ( .A1(n8036), .A2(rEIP[13]), .Y(n8062) );
  NAND2X0_RVT U7411 ( .A1(n8064), .A2(n8065), .Y(n7964) );
  NAND2X0_RVT U7412 ( .A1(n8035), .A2(rEIP[13]), .Y(n8065) );
  NAND2X0_RVT U7413 ( .A1(n8036), .A2(rEIP[14]), .Y(n8064) );
  NAND2X0_RVT U7414 ( .A1(n8066), .A2(n8067), .Y(n7967) );
  NAND2X0_RVT U7415 ( .A1(n8035), .A2(rEIP[14]), .Y(n8067) );
  NAND2X0_RVT U7416 ( .A1(n8036), .A2(rEIP[15]), .Y(n8066) );
  NAND2X0_RVT U7417 ( .A1(n8068), .A2(n8069), .Y(n7972) );
  NAND2X0_RVT U7418 ( .A1(n8035), .A2(rEIP[15]), .Y(n8069) );
  NAND2X0_RVT U7419 ( .A1(n8036), .A2(rEIP[16]), .Y(n8068) );
  NAND2X0_RVT U7420 ( .A1(n8070), .A2(n8071), .Y(n7975) );
  NAND2X0_RVT U7421 ( .A1(n8035), .A2(rEIP[16]), .Y(n8071) );
  NAND2X0_RVT U7422 ( .A1(n8036), .A2(rEIP[17]), .Y(n8070) );
  NAND2X0_RVT U7423 ( .A1(n8072), .A2(n8073), .Y(n7980) );
  NAND2X0_RVT U7424 ( .A1(n8035), .A2(rEIP[17]), .Y(n8073) );
  NAND2X0_RVT U7425 ( .A1(n8036), .A2(rEIP[18]), .Y(n8072) );
  NAND2X0_RVT U7426 ( .A1(n8074), .A2(n8075), .Y(n7983) );
  NAND2X0_RVT U7427 ( .A1(n8035), .A2(rEIP[18]), .Y(n8075) );
  NAND2X0_RVT U7428 ( .A1(n8036), .A2(rEIP[19]), .Y(n8074) );
  NAND2X0_RVT U7429 ( .A1(n8076), .A2(n8077), .Y(n7988) );
  NAND2X0_RVT U7430 ( .A1(n8035), .A2(rEIP[19]), .Y(n8077) );
  NAND2X0_RVT U7431 ( .A1(n8036), .A2(rEIP[20]), .Y(n8076) );
  NAND2X0_RVT U7432 ( .A1(n8078), .A2(n8079), .Y(n7991) );
  NAND2X0_RVT U7433 ( .A1(n8035), .A2(rEIP[20]), .Y(n8079) );
  NAND2X0_RVT U7434 ( .A1(n8036), .A2(rEIP[21]), .Y(n8078) );
  NAND2X0_RVT U7435 ( .A1(n8080), .A2(n8081), .Y(n7996) );
  NAND2X0_RVT U7436 ( .A1(n8035), .A2(rEIP[21]), .Y(n8081) );
  NAND2X0_RVT U7437 ( .A1(n8036), .A2(rEIP[22]), .Y(n8080) );
  NAND2X0_RVT U7438 ( .A1(n8082), .A2(n8083), .Y(n7999) );
  NAND2X0_RVT U7439 ( .A1(n8035), .A2(rEIP[22]), .Y(n8083) );
  NAND2X0_RVT U7440 ( .A1(n8036), .A2(rEIP[23]), .Y(n8082) );
  NAND2X0_RVT U7441 ( .A1(n8084), .A2(n8085), .Y(n8004) );
  NAND2X0_RVT U7442 ( .A1(n8035), .A2(rEIP[23]), .Y(n8085) );
  NAND2X0_RVT U7443 ( .A1(n8036), .A2(rEIP[24]), .Y(n8084) );
  NAND2X0_RVT U7444 ( .A1(n8086), .A2(n8087), .Y(n8007) );
  NAND2X0_RVT U7445 ( .A1(n8035), .A2(rEIP[24]), .Y(n8087) );
  NAND2X0_RVT U7446 ( .A1(n8036), .A2(rEIP[25]), .Y(n8086) );
  NAND2X0_RVT U7447 ( .A1(n8088), .A2(n8089), .Y(n8012) );
  NAND2X0_RVT U7448 ( .A1(n8035), .A2(rEIP[25]), .Y(n8089) );
  NAND2X0_RVT U7449 ( .A1(n8036), .A2(rEIP[26]), .Y(n8088) );
  NAND2X0_RVT U7450 ( .A1(n8090), .A2(n8091), .Y(n8015) );
  NAND2X0_RVT U7451 ( .A1(n8035), .A2(rEIP[26]), .Y(n8091) );
  NAND2X0_RVT U7452 ( .A1(n8036), .A2(rEIP[27]), .Y(n8090) );
  NAND2X0_RVT U7453 ( .A1(n8092), .A2(n8093), .Y(n8020) );
  NAND2X0_RVT U7454 ( .A1(n8035), .A2(rEIP[27]), .Y(n8093) );
  NAND2X0_RVT U7455 ( .A1(n8036), .A2(rEIP[28]), .Y(n8092) );
  NAND2X0_RVT U7456 ( .A1(n8094), .A2(n8095), .Y(n8023) );
  NAND2X0_RVT U7457 ( .A1(n8035), .A2(rEIP[28]), .Y(n8095) );
  NAND2X0_RVT U7458 ( .A1(n8036), .A2(rEIP[29]), .Y(n8094) );
  NAND2X0_RVT U7459 ( .A1(n8096), .A2(n8097), .Y(n8031) );
  NAND2X0_RVT U7460 ( .A1(n8035), .A2(rEIP[30]), .Y(n8097) );
  NAND2X0_RVT U7461 ( .A1(n8036), .A2(rEIP[31]), .Y(n8096) );
  NAND2X0_RVT U7462 ( .A1(n5276), .A2(Address[29]), .Y(n8029) );
  NAND4X0_RVT U7463 ( .A1(n6539), .A2(n8098), .A3(n8099), .A4(n8100), .Y(n4558) );
  NAND2X0_RVT U7464 ( .A1(n7213), .A2(n5479), .Y(n8100) );
  NAND4X0_RVT U7465 ( .A1(n8101), .A2(n8102), .A3(n8103), .A4(n8104), .Y(n7213) );
  NAND2X0_RVT U7466 ( .A1(n8105), .A2(n5118), .Y(n8104) );
  NAND2X0_RVT U7467 ( .A1(n8106), .A2(n8107), .Y(n8103) );
  NAND2X0_RVT U7468 ( .A1(n8108), .A2(n5055), .Y(n8102) );
  NAND2X0_RVT U7469 ( .A1(rEIP[0]), .A2(n8109), .Y(n8101) );
  NAND2X0_RVT U7470 ( .A1(n8110), .A2(n6544), .Y(n8099) );
  XOR2X1_RVT U7471 ( .A1(n8111), .A2(n6543), .Y(n6544) );
  OR2X1_RVT U7472 ( .A1(n8107), .A2(n8112), .Y(n8111) );
  NAND2X0_RVT U7473 ( .A1(n8113), .A2(n5055), .Y(n8098) );
  NAND2X0_RVT U7474 ( .A1(rEIP[0]), .A2(n8114), .Y(n6539) );
  NAND4X0_RVT U7475 ( .A1(n6720), .A2(n8115), .A3(n8116), .A4(n8117), .Y(n4557) );
  NAND2X0_RVT U7476 ( .A1(n7232), .A2(n5479), .Y(n8117) );
  XOR2X1_RVT U7477 ( .A1(n8118), .A2(n8119), .Y(n7232) );
  NAND2X0_RVT U7478 ( .A1(n8110), .A2(n6729), .Y(n8116) );
  XOR3X1_RVT U7479 ( .A1(n8120), .A2(n8121), .A3(n6724), .Y(n6729) );
  NAND2X0_RVT U7480 ( .A1(n8113), .A2(n5063), .Y(n8115) );
  NAND2X0_RVT U7481 ( .A1(rEIP[1]), .A2(n8114), .Y(n6720) );
  NAND4X0_RVT U7482 ( .A1(n6714), .A2(n8122), .A3(n8123), .A4(n8124), .Y(n4556) );
  NAND2X0_RVT U7483 ( .A1(n7248), .A2(n5479), .Y(n8124) );
  XOR3X1_RVT U7484 ( .A1(n8125), .A2(n8126), .A3(n8127), .Y(n7248) );
  NAND2X0_RVT U7485 ( .A1(n8110), .A2(n6719), .Y(n8123) );
  XOR3X1_RVT U7486 ( .A1(n8128), .A2(n8129), .A3(n6718), .Y(n6719) );
  NAND2X0_RVT U7487 ( .A1(n8113), .A2(n5062), .Y(n8122) );
  NAND2X0_RVT U7488 ( .A1(rEIP[2]), .A2(n8114), .Y(n6714) );
  NAND4X0_RVT U7489 ( .A1(n6708), .A2(n8130), .A3(n8131), .A4(n8132), .Y(n4555) );
  NAND2X0_RVT U7490 ( .A1(n7281), .A2(n5479), .Y(n8132) );
  NAND3X0_RVT U7491 ( .A1(n8133), .A2(n8134), .A3(n8135), .Y(n7281) );
  XNOR2X1_RVT U7492 ( .A1(n8136), .A2(n8137), .Y(n8135) );
  NAND2X0_RVT U7493 ( .A1(n8105), .A2(n5119), .Y(n8134) );
  NAND2X0_RVT U7494 ( .A1(n8106), .A2(n8138), .Y(n8133) );
  NAND2X0_RVT U7495 ( .A1(n8110), .A2(n6713), .Y(n8131) );
  XOR3X1_RVT U7496 ( .A1(n8139), .A2(n8140), .A3(n6712), .Y(n6713) );
  NAND2X0_RVT U7497 ( .A1(n8113), .A2(n5061), .Y(n8130) );
  NAND2X0_RVT U7498 ( .A1(rEIP[3]), .A2(n8114), .Y(n6708) );
  NAND4X0_RVT U7499 ( .A1(n6702), .A2(n8141), .A3(n8142), .A4(n8143), .Y(n4554) );
  NAND2X0_RVT U7500 ( .A1(n7292), .A2(n5479), .Y(n8143) );
  NAND3X0_RVT U7501 ( .A1(n8144), .A2(n8145), .A3(n8146), .Y(n7292) );
  XNOR2X1_RVT U7502 ( .A1(n8147), .A2(n8148), .Y(n8146) );
  NAND2X0_RVT U7503 ( .A1(n8105), .A2(n5120), .Y(n8145) );
  NAND2X0_RVT U7504 ( .A1(n8106), .A2(n8149), .Y(n8144) );
  NAND2X0_RVT U7505 ( .A1(n8110), .A2(n6707), .Y(n8142) );
  XOR3X1_RVT U7506 ( .A1(n8150), .A2(n8151), .A3(n6706), .Y(n6707) );
  NAND2X0_RVT U7507 ( .A1(n8113), .A2(n5060), .Y(n8141) );
  NAND2X0_RVT U7508 ( .A1(rEIP[4]), .A2(n8114), .Y(n6702) );
  NAND4X0_RVT U7509 ( .A1(n6696), .A2(n8152), .A3(n8153), .A4(n8154), .Y(n4553) );
  NAND2X0_RVT U7510 ( .A1(n7303), .A2(n5479), .Y(n8154) );
  NAND3X0_RVT U7511 ( .A1(n8155), .A2(n8156), .A3(n8157), .Y(n7303) );
  XNOR2X1_RVT U7512 ( .A1(n8158), .A2(n8159), .Y(n8157) );
  NAND2X0_RVT U7513 ( .A1(n8105), .A2(n5121), .Y(n8156) );
  NAND2X0_RVT U7514 ( .A1(n8106), .A2(n8160), .Y(n8155) );
  NAND2X0_RVT U7515 ( .A1(n8110), .A2(n6701), .Y(n8153) );
  XOR3X1_RVT U7516 ( .A1(n8161), .A2(n8162), .A3(n6700), .Y(n6701) );
  NAND2X0_RVT U7517 ( .A1(n8113), .A2(n5059), .Y(n8152) );
  NAND2X0_RVT U7518 ( .A1(rEIP[5]), .A2(n8114), .Y(n6696) );
  NAND4X0_RVT U7519 ( .A1(n6690), .A2(n8163), .A3(n8164), .A4(n8165), .Y(n4552) );
  NAND2X0_RVT U7520 ( .A1(n7314), .A2(n5479), .Y(n8165) );
  NAND3X0_RVT U7521 ( .A1(n8166), .A2(n8167), .A3(n8168), .Y(n7314) );
  XNOR2X1_RVT U7522 ( .A1(n8169), .A2(n8170), .Y(n8168) );
  NAND2X0_RVT U7523 ( .A1(n8105), .A2(n5122), .Y(n8167) );
  NAND2X0_RVT U7524 ( .A1(n8106), .A2(n8171), .Y(n8166) );
  NAND2X0_RVT U7525 ( .A1(n8110), .A2(n6695), .Y(n8164) );
  XOR3X1_RVT U7526 ( .A1(n8172), .A2(n8173), .A3(n6694), .Y(n6695) );
  NAND2X0_RVT U7527 ( .A1(n8113), .A2(n5058), .Y(n8163) );
  NAND2X0_RVT U7528 ( .A1(rEIP[6]), .A2(n8114), .Y(n6690) );
  NAND4X0_RVT U7529 ( .A1(n6684), .A2(n8174), .A3(n8175), .A4(n8176), .Y(n4551) );
  NAND2X0_RVT U7530 ( .A1(n7325), .A2(n5479), .Y(n8176) );
  NAND3X0_RVT U7531 ( .A1(n8177), .A2(n8178), .A3(n8179), .Y(n7325) );
  XNOR2X1_RVT U7532 ( .A1(n8180), .A2(n8181), .Y(n8179) );
  NAND2X0_RVT U7533 ( .A1(n8105), .A2(n5049), .Y(n8178) );
  NAND2X0_RVT U7534 ( .A1(n8106), .A2(n8182), .Y(n8177) );
  NAND2X0_RVT U7535 ( .A1(n8110), .A2(n6689), .Y(n8175) );
  XNOR3X1_RVT U7536 ( .A1(n8183), .A2(n8184), .A3(n8185), .Y(n6689) );
  NAND2X0_RVT U7537 ( .A1(n8113), .A2(n5057), .Y(n8174) );
  NAND2X0_RVT U7538 ( .A1(rEIP[7]), .A2(n8114), .Y(n6684) );
  NAND4X0_RVT U7539 ( .A1(n6678), .A2(n8186), .A3(n8187), .A4(n8188), .Y(n4550) );
  NAND2X0_RVT U7540 ( .A1(n7336), .A2(n5479), .Y(n8188) );
  XOR2X1_RVT U7541 ( .A1(n8189), .A2(n8190), .Y(n7336) );
  NAND2X0_RVT U7542 ( .A1(n8110), .A2(n6683), .Y(n8187) );
  XNOR3X1_RVT U7543 ( .A1(n8191), .A2(n8192), .A3(n6682), .Y(n6683) );
  NAND2X0_RVT U7544 ( .A1(n8113), .A2(n5064), .Y(n8186) );
  NAND2X0_RVT U7545 ( .A1(rEIP[8]), .A2(n8114), .Y(n6678) );
  NAND4X0_RVT U7546 ( .A1(n6672), .A2(n8193), .A3(n8194), .A4(n8195), .Y(n4549) );
  NAND2X0_RVT U7547 ( .A1(n7347), .A2(n5479), .Y(n8195) );
  XNOR2X1_RVT U7548 ( .A1(n8196), .A2(n8197), .Y(n7347) );
  NAND2X0_RVT U7549 ( .A1(n8189), .A2(n8190), .Y(n8196) );
  NAND2X0_RVT U7550 ( .A1(n8110), .A2(n6677), .Y(n8194) );
  XNOR3X1_RVT U7551 ( .A1(n8192), .A2(n6676), .A3(n8198), .Y(n6677) );
  NAND2X0_RVT U7552 ( .A1(n8113), .A2(n5065), .Y(n8193) );
  NAND2X0_RVT U7553 ( .A1(rEIP[9]), .A2(n8114), .Y(n6672) );
  NAND4X0_RVT U7554 ( .A1(n6666), .A2(n8199), .A3(n8200), .A4(n8201), .Y(n4548) );
  NAND2X0_RVT U7555 ( .A1(n7358), .A2(n5479), .Y(n8201) );
  XOR2X1_RVT U7556 ( .A1(n8202), .A2(n8203), .Y(n7358) );
  NAND2X0_RVT U7557 ( .A1(n8110), .A2(n6671), .Y(n8200) );
  XNOR3X1_RVT U7558 ( .A1(n8192), .A2(n6670), .A3(n8204), .Y(n6671) );
  NAND2X0_RVT U7559 ( .A1(n8113), .A2(n5066), .Y(n8199) );
  NAND2X0_RVT U7560 ( .A1(rEIP[10]), .A2(n8114), .Y(n6666) );
  NAND4X0_RVT U7561 ( .A1(n6660), .A2(n8205), .A3(n8206), .A4(n8207), .Y(n4547) );
  NAND2X0_RVT U7562 ( .A1(n7369), .A2(n5479), .Y(n8207) );
  XNOR2X1_RVT U7563 ( .A1(n8208), .A2(n8209), .Y(n7369) );
  NAND2X0_RVT U7564 ( .A1(n8202), .A2(n8203), .Y(n8208) );
  NAND2X0_RVT U7565 ( .A1(n8110), .A2(n6665), .Y(n8206) );
  XNOR3X1_RVT U7566 ( .A1(n8192), .A2(n6664), .A3(n8210), .Y(n6665) );
  NAND2X0_RVT U7567 ( .A1(n8113), .A2(n5067), .Y(n8205) );
  NAND2X0_RVT U7568 ( .A1(rEIP[11]), .A2(n8114), .Y(n6660) );
  NAND4X0_RVT U7569 ( .A1(n6654), .A2(n8211), .A3(n8212), .A4(n8213), .Y(n4546) );
  NAND2X0_RVT U7570 ( .A1(n7380), .A2(n5479), .Y(n8213) );
  XOR2X1_RVT U7571 ( .A1(n8214), .A2(n8215), .Y(n7380) );
  NAND2X0_RVT U7572 ( .A1(n8110), .A2(n6659), .Y(n8212) );
  XNOR3X1_RVT U7573 ( .A1(n8192), .A2(n6658), .A3(n8216), .Y(n6659) );
  NAND2X0_RVT U7574 ( .A1(n8113), .A2(n5068), .Y(n8211) );
  NAND2X0_RVT U7575 ( .A1(rEIP[12]), .A2(n8114), .Y(n6654) );
  NAND4X0_RVT U7576 ( .A1(n6648), .A2(n8217), .A3(n8218), .A4(n8219), .Y(n4545) );
  NAND2X0_RVT U7577 ( .A1(n7391), .A2(n5479), .Y(n8219) );
  XNOR2X1_RVT U7578 ( .A1(n8220), .A2(n8221), .Y(n7391) );
  NAND2X0_RVT U7579 ( .A1(n8214), .A2(n8215), .Y(n8220) );
  NAND2X0_RVT U7580 ( .A1(n8110), .A2(n6653), .Y(n8218) );
  XNOR3X1_RVT U7581 ( .A1(n8192), .A2(n6652), .A3(n8222), .Y(n6653) );
  NAND2X0_RVT U7582 ( .A1(n8113), .A2(n5069), .Y(n8217) );
  NAND2X0_RVT U7583 ( .A1(rEIP[13]), .A2(n8114), .Y(n6648) );
  NAND4X0_RVT U7584 ( .A1(n6642), .A2(n8223), .A3(n8224), .A4(n8225), .Y(n4544) );
  NAND2X0_RVT U7585 ( .A1(n7402), .A2(n5479), .Y(n8225) );
  XOR2X1_RVT U7586 ( .A1(n8226), .A2(n8227), .Y(n7402) );
  NAND2X0_RVT U7587 ( .A1(n8110), .A2(n6647), .Y(n8224) );
  XNOR3X1_RVT U7588 ( .A1(n8192), .A2(n6646), .A3(n8228), .Y(n6647) );
  NAND2X0_RVT U7589 ( .A1(n8113), .A2(n5070), .Y(n8223) );
  NAND2X0_RVT U7590 ( .A1(rEIP[14]), .A2(n8114), .Y(n6642) );
  NAND4X0_RVT U7591 ( .A1(n6636), .A2(n8229), .A3(n8230), .A4(n8231), .Y(n4543) );
  NAND2X0_RVT U7592 ( .A1(n7413), .A2(n5479), .Y(n8231) );
  XNOR2X1_RVT U7593 ( .A1(n8232), .A2(n8233), .Y(n7413) );
  NAND2X0_RVT U7594 ( .A1(n8226), .A2(n8227), .Y(n8232) );
  NAND2X0_RVT U7595 ( .A1(n8110), .A2(n6641), .Y(n8230) );
  XNOR3X1_RVT U7596 ( .A1(n8192), .A2(n6640), .A3(n8234), .Y(n6641) );
  NAND2X0_RVT U7597 ( .A1(n8113), .A2(n5071), .Y(n8229) );
  NAND2X0_RVT U7598 ( .A1(rEIP[15]), .A2(n8114), .Y(n6636) );
  NAND4X0_RVT U7599 ( .A1(n6630), .A2(n8235), .A3(n8236), .A4(n8237), .Y(n4542) );
  NAND2X0_RVT U7600 ( .A1(n7424), .A2(n5479), .Y(n8237) );
  XOR2X1_RVT U7601 ( .A1(n8238), .A2(n8239), .Y(n7424) );
  NAND2X0_RVT U7602 ( .A1(n8110), .A2(n6635), .Y(n8236) );
  XNOR3X1_RVT U7603 ( .A1(n8192), .A2(n6634), .A3(n8240), .Y(n6635) );
  NAND2X0_RVT U7604 ( .A1(n8113), .A2(n5072), .Y(n8235) );
  NAND2X0_RVT U7605 ( .A1(rEIP[16]), .A2(n8114), .Y(n6630) );
  NAND4X0_RVT U7606 ( .A1(n6624), .A2(n8241), .A3(n8242), .A4(n8243), .Y(n4541) );
  NAND2X0_RVT U7607 ( .A1(n7441), .A2(n5479), .Y(n8243) );
  XNOR2X1_RVT U7608 ( .A1(n8244), .A2(n8245), .Y(n7441) );
  NAND2X0_RVT U7609 ( .A1(n8238), .A2(n8239), .Y(n8244) );
  NAND2X0_RVT U7610 ( .A1(n8110), .A2(n6629), .Y(n8242) );
  XNOR3X1_RVT U7611 ( .A1(n8192), .A2(n6628), .A3(n8246), .Y(n6629) );
  NAND2X0_RVT U7612 ( .A1(n8113), .A2(n5073), .Y(n8241) );
  NAND2X0_RVT U7613 ( .A1(rEIP[17]), .A2(n8114), .Y(n6624) );
  NAND4X0_RVT U7614 ( .A1(n6618), .A2(n8247), .A3(n8248), .A4(n8249), .Y(n4540) );
  NAND2X0_RVT U7615 ( .A1(n7457), .A2(n5479), .Y(n8249) );
  XOR2X1_RVT U7616 ( .A1(n8250), .A2(n8251), .Y(n7457) );
  NAND2X0_RVT U7617 ( .A1(n8110), .A2(n6623), .Y(n8248) );
  XNOR3X1_RVT U7618 ( .A1(n8192), .A2(n6622), .A3(n8252), .Y(n6623) );
  NAND2X0_RVT U7619 ( .A1(n8113), .A2(n5074), .Y(n8247) );
  NAND2X0_RVT U7620 ( .A1(rEIP[18]), .A2(n8114), .Y(n6618) );
  NAND4X0_RVT U7621 ( .A1(n6612), .A2(n8253), .A3(n8254), .A4(n8255), .Y(n4539) );
  NAND2X0_RVT U7622 ( .A1(n7473), .A2(n5479), .Y(n8255) );
  XNOR2X1_RVT U7623 ( .A1(n8256), .A2(n8257), .Y(n7473) );
  NAND2X0_RVT U7624 ( .A1(n8250), .A2(n8251), .Y(n8256) );
  NAND2X0_RVT U7625 ( .A1(n8110), .A2(n6617), .Y(n8254) );
  XNOR3X1_RVT U7626 ( .A1(n8192), .A2(n6616), .A3(n8258), .Y(n6617) );
  NAND2X0_RVT U7627 ( .A1(n8113), .A2(n5075), .Y(n8253) );
  NAND2X0_RVT U7628 ( .A1(rEIP[19]), .A2(n8114), .Y(n6612) );
  NAND4X0_RVT U7629 ( .A1(n6606), .A2(n8259), .A3(n8260), .A4(n8261), .Y(n4538) );
  NAND2X0_RVT U7630 ( .A1(n7488), .A2(n5479), .Y(n8261) );
  XOR2X1_RVT U7631 ( .A1(n8262), .A2(n8263), .Y(n7488) );
  NAND2X0_RVT U7632 ( .A1(n8110), .A2(n6611), .Y(n8260) );
  XNOR3X1_RVT U7633 ( .A1(n8192), .A2(n6610), .A3(n8264), .Y(n6611) );
  NAND2X0_RVT U7634 ( .A1(n8113), .A2(n5076), .Y(n8259) );
  NAND2X0_RVT U7635 ( .A1(rEIP[20]), .A2(n8114), .Y(n6606) );
  NAND4X0_RVT U7636 ( .A1(n6600), .A2(n8265), .A3(n8266), .A4(n8267), .Y(n4537) );
  NAND2X0_RVT U7637 ( .A1(n7504), .A2(n5479), .Y(n8267) );
  XNOR2X1_RVT U7638 ( .A1(n8268), .A2(n8269), .Y(n7504) );
  NAND2X0_RVT U7639 ( .A1(n8262), .A2(n8263), .Y(n8268) );
  NAND2X0_RVT U7640 ( .A1(n8110), .A2(n6605), .Y(n8266) );
  XNOR3X1_RVT U7641 ( .A1(n8192), .A2(n6604), .A3(n8270), .Y(n6605) );
  NAND2X0_RVT U7642 ( .A1(n8113), .A2(n5077), .Y(n8265) );
  NAND2X0_RVT U7643 ( .A1(rEIP[21]), .A2(n8114), .Y(n6600) );
  NAND4X0_RVT U7644 ( .A1(n6594), .A2(n8271), .A3(n8272), .A4(n8273), .Y(n4536) );
  NAND2X0_RVT U7645 ( .A1(n7520), .A2(n5479), .Y(n8273) );
  XOR2X1_RVT U7646 ( .A1(n8274), .A2(n8275), .Y(n7520) );
  NAND2X0_RVT U7647 ( .A1(n8110), .A2(n6599), .Y(n8272) );
  XNOR3X1_RVT U7648 ( .A1(n8192), .A2(n6598), .A3(n8276), .Y(n6599) );
  NAND2X0_RVT U7649 ( .A1(n8113), .A2(n5078), .Y(n8271) );
  NAND2X0_RVT U7650 ( .A1(rEIP[22]), .A2(n8114), .Y(n6594) );
  NAND4X0_RVT U7651 ( .A1(n6588), .A2(n8277), .A3(n8278), .A4(n8279), .Y(n4535) );
  NAND2X0_RVT U7652 ( .A1(n7536), .A2(n5479), .Y(n8279) );
  XNOR2X1_RVT U7653 ( .A1(n8280), .A2(n8281), .Y(n7536) );
  NAND2X0_RVT U7654 ( .A1(n8274), .A2(n8275), .Y(n8280) );
  NAND2X0_RVT U7655 ( .A1(n8110), .A2(n6593), .Y(n8278) );
  XNOR3X1_RVT U7656 ( .A1(n8192), .A2(n6592), .A3(n8282), .Y(n6593) );
  NAND2X0_RVT U7657 ( .A1(n8113), .A2(n5079), .Y(n8277) );
  NAND2X0_RVT U7658 ( .A1(rEIP[23]), .A2(n8114), .Y(n6588) );
  NAND4X0_RVT U7659 ( .A1(n6582), .A2(n8283), .A3(n8284), .A4(n8285), .Y(n4534) );
  NAND2X0_RVT U7660 ( .A1(n7553), .A2(n5479), .Y(n8285) );
  XOR2X1_RVT U7661 ( .A1(n8286), .A2(n8287), .Y(n7553) );
  NAND2X0_RVT U7662 ( .A1(n8110), .A2(n6587), .Y(n8284) );
  XNOR3X1_RVT U7663 ( .A1(n8192), .A2(n6586), .A3(n8288), .Y(n6587) );
  NAND2X0_RVT U7664 ( .A1(n8113), .A2(n5080), .Y(n8283) );
  NAND2X0_RVT U7665 ( .A1(rEIP[24]), .A2(n8114), .Y(n6582) );
  NAND4X0_RVT U7666 ( .A1(n6576), .A2(n8289), .A3(n8290), .A4(n8291), .Y(n4533) );
  NAND2X0_RVT U7667 ( .A1(n7571), .A2(n5479), .Y(n8291) );
  XNOR2X1_RVT U7668 ( .A1(n8292), .A2(n8293), .Y(n7571) );
  NAND2X0_RVT U7669 ( .A1(n8286), .A2(n8287), .Y(n8292) );
  NAND2X0_RVT U7670 ( .A1(n8110), .A2(n6581), .Y(n8290) );
  XNOR3X1_RVT U7671 ( .A1(n8192), .A2(n6580), .A3(n8294), .Y(n6581) );
  NAND2X0_RVT U7672 ( .A1(n8113), .A2(n5081), .Y(n8289) );
  NAND2X0_RVT U7673 ( .A1(rEIP[25]), .A2(n8114), .Y(n6576) );
  NAND4X0_RVT U7674 ( .A1(n6570), .A2(n8295), .A3(n8296), .A4(n8297), .Y(n4532) );
  NAND2X0_RVT U7675 ( .A1(n7589), .A2(n5479), .Y(n8297) );
  XOR2X1_RVT U7676 ( .A1(n8298), .A2(n8299), .Y(n7589) );
  NAND2X0_RVT U7677 ( .A1(n8110), .A2(n6575), .Y(n8296) );
  XNOR3X1_RVT U7678 ( .A1(n8192), .A2(n6574), .A3(n8300), .Y(n6575) );
  NAND2X0_RVT U7679 ( .A1(n8113), .A2(n5082), .Y(n8295) );
  NAND2X0_RVT U7680 ( .A1(rEIP[26]), .A2(n8114), .Y(n6570) );
  NAND4X0_RVT U7681 ( .A1(n6564), .A2(n8301), .A3(n8302), .A4(n8303), .Y(n4531) );
  NAND2X0_RVT U7682 ( .A1(n7607), .A2(n5479), .Y(n8303) );
  XNOR2X1_RVT U7683 ( .A1(n8304), .A2(n8305), .Y(n7607) );
  NAND2X0_RVT U7684 ( .A1(n8298), .A2(n8299), .Y(n8304) );
  NAND2X0_RVT U7685 ( .A1(n8110), .A2(n6569), .Y(n8302) );
  XNOR3X1_RVT U7686 ( .A1(n8192), .A2(n6568), .A3(n8306), .Y(n6569) );
  NAND2X0_RVT U7687 ( .A1(n8113), .A2(n5083), .Y(n8301) );
  NAND2X0_RVT U7688 ( .A1(rEIP[27]), .A2(n8114), .Y(n6564) );
  NAND4X0_RVT U7689 ( .A1(n6558), .A2(n8307), .A3(n8308), .A4(n8309), .Y(n4530) );
  NAND2X0_RVT U7690 ( .A1(n7625), .A2(n5479), .Y(n8309) );
  XOR2X1_RVT U7691 ( .A1(n8310), .A2(n8311), .Y(n7625) );
  NAND2X0_RVT U7692 ( .A1(n8110), .A2(n6563), .Y(n8308) );
  XNOR3X1_RVT U7693 ( .A1(n8192), .A2(n6562), .A3(n8312), .Y(n6563) );
  NAND2X0_RVT U7694 ( .A1(n8113), .A2(n5084), .Y(n8307) );
  NAND2X0_RVT U7695 ( .A1(rEIP[28]), .A2(n8114), .Y(n6558) );
  NAND4X0_RVT U7696 ( .A1(n6552), .A2(n8313), .A3(n8314), .A4(n8315), .Y(n4529) );
  NAND2X0_RVT U7697 ( .A1(n7643), .A2(n5479), .Y(n8315) );
  XNOR2X1_RVT U7698 ( .A1(n8316), .A2(n8317), .Y(n7643) );
  NAND2X0_RVT U7699 ( .A1(n8310), .A2(n8311), .Y(n8316) );
  NAND2X0_RVT U7700 ( .A1(n8110), .A2(n6557), .Y(n8314) );
  XNOR3X1_RVT U7701 ( .A1(n8192), .A2(n6556), .A3(n8318), .Y(n6557) );
  NAND2X0_RVT U7702 ( .A1(n8113), .A2(n5085), .Y(n8313) );
  NAND2X0_RVT U7703 ( .A1(rEIP[29]), .A2(n8114), .Y(n6552) );
  NAND4X0_RVT U7704 ( .A1(n6546), .A2(n8319), .A3(n8320), .A4(n8321), .Y(n4528) );
  NAND2X0_RVT U7705 ( .A1(n7661), .A2(n5479), .Y(n8321) );
  XOR2X1_RVT U7706 ( .A1(n8322), .A2(n8323), .Y(n7661) );
  NAND2X0_RVT U7707 ( .A1(n8110), .A2(n6551), .Y(n8320) );
  XNOR3X1_RVT U7708 ( .A1(n8192), .A2(n6550), .A3(n8324), .Y(n6551) );
  NAND2X0_RVT U7709 ( .A1(n8113), .A2(n5056), .Y(n8319) );
  NAND2X0_RVT U7710 ( .A1(rEIP[30]), .A2(n8114), .Y(n6546) );
  NAND4X0_RVT U7711 ( .A1(n5315), .A2(n8325), .A3(n8326), .A4(n8327), .Y(n4527) );
  NAND2X0_RVT U7712 ( .A1(n8110), .A2(n5322), .Y(n8327) );
  XNOR3X1_RVT U7713 ( .A1(n8192), .A2(n5320), .A3(n8328), .Y(n5322) );
  NAND2X0_RVT U7714 ( .A1(n8329), .A2(n8330), .Y(n8328) );
  NAND2X0_RVT U7715 ( .A1(n8112), .A2(n8331), .Y(n8330) );
  OR2X1_RVT U7716 ( .A1(n8324), .A2(n6550), .Y(n8331) );
  NAND2X0_RVT U7717 ( .A1(n6550), .A2(n8324), .Y(n8329) );
  NAND2X0_RVT U7718 ( .A1(n8332), .A2(n8333), .Y(n8324) );
  NAND2X0_RVT U7719 ( .A1(n8112), .A2(n8334), .Y(n8333) );
  OR2X1_RVT U7720 ( .A1(n8318), .A2(n6556), .Y(n8334) );
  NAND2X0_RVT U7721 ( .A1(n6556), .A2(n8318), .Y(n8332) );
  NAND2X0_RVT U7722 ( .A1(n8335), .A2(n8336), .Y(n8318) );
  NAND2X0_RVT U7723 ( .A1(n8112), .A2(n8337), .Y(n8336) );
  OR2X1_RVT U7724 ( .A1(n8312), .A2(n6562), .Y(n8337) );
  NAND2X0_RVT U7725 ( .A1(n6562), .A2(n8312), .Y(n8335) );
  NAND2X0_RVT U7726 ( .A1(n8338), .A2(n8339), .Y(n8312) );
  NAND2X0_RVT U7727 ( .A1(n8112), .A2(n8340), .Y(n8339) );
  OR2X1_RVT U7728 ( .A1(n8306), .A2(n6568), .Y(n8340) );
  NAND2X0_RVT U7729 ( .A1(n6568), .A2(n8306), .Y(n8338) );
  NAND2X0_RVT U7730 ( .A1(n8341), .A2(n8342), .Y(n8306) );
  NAND2X0_RVT U7731 ( .A1(n8112), .A2(n8343), .Y(n8342) );
  OR2X1_RVT U7732 ( .A1(n8300), .A2(n6574), .Y(n8343) );
  NAND2X0_RVT U7733 ( .A1(n6574), .A2(n8300), .Y(n8341) );
  NAND2X0_RVT U7734 ( .A1(n8344), .A2(n8345), .Y(n8300) );
  NAND2X0_RVT U7735 ( .A1(n8112), .A2(n8346), .Y(n8345) );
  OR2X1_RVT U7736 ( .A1(n8294), .A2(n6580), .Y(n8346) );
  NAND2X0_RVT U7737 ( .A1(n6580), .A2(n8294), .Y(n8344) );
  NAND2X0_RVT U7738 ( .A1(n8347), .A2(n8348), .Y(n8294) );
  NAND2X0_RVT U7739 ( .A1(n8112), .A2(n8349), .Y(n8348) );
  OR2X1_RVT U7740 ( .A1(n8288), .A2(n6586), .Y(n8349) );
  NAND2X0_RVT U7741 ( .A1(n6586), .A2(n8288), .Y(n8347) );
  NAND2X0_RVT U7742 ( .A1(n8350), .A2(n8351), .Y(n8288) );
  NAND2X0_RVT U7743 ( .A1(n8112), .A2(n8352), .Y(n8351) );
  OR2X1_RVT U7744 ( .A1(n8282), .A2(n6592), .Y(n8352) );
  NAND2X0_RVT U7745 ( .A1(n6592), .A2(n8282), .Y(n8350) );
  NAND2X0_RVT U7746 ( .A1(n8353), .A2(n8354), .Y(n8282) );
  NAND2X0_RVT U7747 ( .A1(n8112), .A2(n8355), .Y(n8354) );
  OR2X1_RVT U7748 ( .A1(n8276), .A2(n6598), .Y(n8355) );
  NAND2X0_RVT U7749 ( .A1(n6598), .A2(n8276), .Y(n8353) );
  NAND2X0_RVT U7750 ( .A1(n8356), .A2(n8357), .Y(n8276) );
  NAND2X0_RVT U7751 ( .A1(n8112), .A2(n8358), .Y(n8357) );
  OR2X1_RVT U7752 ( .A1(n8270), .A2(n6604), .Y(n8358) );
  NAND2X0_RVT U7753 ( .A1(n6604), .A2(n8270), .Y(n8356) );
  NAND2X0_RVT U7754 ( .A1(n8359), .A2(n8360), .Y(n8270) );
  NAND2X0_RVT U7755 ( .A1(n8112), .A2(n8361), .Y(n8360) );
  OR2X1_RVT U7756 ( .A1(n8264), .A2(n6610), .Y(n8361) );
  NAND2X0_RVT U7757 ( .A1(n6610), .A2(n8264), .Y(n8359) );
  NAND2X0_RVT U7758 ( .A1(n8362), .A2(n8363), .Y(n8264) );
  NAND2X0_RVT U7759 ( .A1(n8112), .A2(n8364), .Y(n8363) );
  OR2X1_RVT U7760 ( .A1(n8258), .A2(n6616), .Y(n8364) );
  NAND2X0_RVT U7761 ( .A1(n6616), .A2(n8258), .Y(n8362) );
  NAND2X0_RVT U7762 ( .A1(n8365), .A2(n8366), .Y(n8258) );
  NAND2X0_RVT U7763 ( .A1(n8112), .A2(n8367), .Y(n8366) );
  OR2X1_RVT U7764 ( .A1(n8252), .A2(n6622), .Y(n8367) );
  NAND2X0_RVT U7765 ( .A1(n6622), .A2(n8252), .Y(n8365) );
  NAND2X0_RVT U7766 ( .A1(n8368), .A2(n8369), .Y(n8252) );
  NAND2X0_RVT U7767 ( .A1(n8112), .A2(n8370), .Y(n8369) );
  OR2X1_RVT U7768 ( .A1(n8246), .A2(n6628), .Y(n8370) );
  NAND2X0_RVT U7769 ( .A1(n6628), .A2(n8246), .Y(n8368) );
  NAND2X0_RVT U7770 ( .A1(n8371), .A2(n8372), .Y(n8246) );
  NAND2X0_RVT U7771 ( .A1(n8112), .A2(n8373), .Y(n8372) );
  OR2X1_RVT U7772 ( .A1(n8240), .A2(n6634), .Y(n8373) );
  NAND2X0_RVT U7773 ( .A1(n6634), .A2(n8240), .Y(n8371) );
  NAND2X0_RVT U7774 ( .A1(n8374), .A2(n8375), .Y(n8240) );
  NAND2X0_RVT U7775 ( .A1(n8112), .A2(n8376), .Y(n8375) );
  OR2X1_RVT U7776 ( .A1(n8234), .A2(n6640), .Y(n8376) );
  NAND2X0_RVT U7777 ( .A1(n6640), .A2(n8234), .Y(n8374) );
  NAND2X0_RVT U7778 ( .A1(n8377), .A2(n8378), .Y(n8234) );
  NAND2X0_RVT U7779 ( .A1(n8112), .A2(n8379), .Y(n8378) );
  OR2X1_RVT U7780 ( .A1(n8228), .A2(n6646), .Y(n8379) );
  NAND2X0_RVT U7781 ( .A1(n6646), .A2(n8228), .Y(n8377) );
  NAND2X0_RVT U7782 ( .A1(n8380), .A2(n8381), .Y(n8228) );
  NAND2X0_RVT U7783 ( .A1(n8112), .A2(n8382), .Y(n8381) );
  OR2X1_RVT U7784 ( .A1(n8222), .A2(n6652), .Y(n8382) );
  NAND2X0_RVT U7785 ( .A1(n6652), .A2(n8222), .Y(n8380) );
  NAND2X0_RVT U7786 ( .A1(n8383), .A2(n8384), .Y(n8222) );
  NAND2X0_RVT U7787 ( .A1(n8112), .A2(n8385), .Y(n8384) );
  OR2X1_RVT U7788 ( .A1(n8216), .A2(n6658), .Y(n8385) );
  NAND2X0_RVT U7789 ( .A1(n6658), .A2(n8216), .Y(n8383) );
  NAND2X0_RVT U7790 ( .A1(n8386), .A2(n8387), .Y(n8216) );
  NAND2X0_RVT U7791 ( .A1(n8112), .A2(n8388), .Y(n8387) );
  OR2X1_RVT U7792 ( .A1(n8210), .A2(n6664), .Y(n8388) );
  NAND2X0_RVT U7793 ( .A1(n6664), .A2(n8210), .Y(n8386) );
  NAND2X0_RVT U7794 ( .A1(n8389), .A2(n8390), .Y(n8210) );
  NAND2X0_RVT U7795 ( .A1(n8112), .A2(n8391), .Y(n8390) );
  OR2X1_RVT U7796 ( .A1(n8204), .A2(n6670), .Y(n8391) );
  NAND2X0_RVT U7797 ( .A1(n6670), .A2(n8204), .Y(n8389) );
  NAND2X0_RVT U7798 ( .A1(n8392), .A2(n8393), .Y(n8204) );
  NAND2X0_RVT U7799 ( .A1(n8112), .A2(n8394), .Y(n8393) );
  OR2X1_RVT U7800 ( .A1(n8198), .A2(n6676), .Y(n8394) );
  NAND2X0_RVT U7801 ( .A1(n6676), .A2(n8198), .Y(n8392) );
  NAND2X0_RVT U7802 ( .A1(n8395), .A2(n8396), .Y(n8198) );
  NAND2X0_RVT U7803 ( .A1(n8112), .A2(n8397), .Y(n8396) );
  OR2X1_RVT U7804 ( .A1(n8191), .A2(n6682), .Y(n8397) );
  NAND2X0_RVT U7805 ( .A1(n6682), .A2(n8191), .Y(n8395) );
  NAND2X0_RVT U7806 ( .A1(n8398), .A2(n8399), .Y(n8191) );
  NAND2X0_RVT U7807 ( .A1(n8184), .A2(n8400), .Y(n8399) );
  OR2X1_RVT U7808 ( .A1(n8183), .A2(n6688), .Y(n8400) );
  AND2X1_RVT U7809 ( .A1(n8401), .A2(n8182), .Y(n8184) );
  NAND2X0_RVT U7810 ( .A1(n6688), .A2(n8183), .Y(n8398) );
  NAND2X0_RVT U7811 ( .A1(n8402), .A2(n8403), .Y(n8183) );
  NAND2X0_RVT U7812 ( .A1(n8173), .A2(n8404), .Y(n8403) );
  OR2X1_RVT U7813 ( .A1(n8172), .A2(n6694), .Y(n8404) );
  AND2X1_RVT U7814 ( .A1(n8401), .A2(n8171), .Y(n8173) );
  NAND2X0_RVT U7815 ( .A1(n6694), .A2(n8172), .Y(n8402) );
  NAND2X0_RVT U7816 ( .A1(n8405), .A2(n8406), .Y(n8172) );
  NAND2X0_RVT U7817 ( .A1(n8162), .A2(n8407), .Y(n8406) );
  OR2X1_RVT U7818 ( .A1(n8161), .A2(n6700), .Y(n8407) );
  AND2X1_RVT U7819 ( .A1(n8401), .A2(n8160), .Y(n8162) );
  NAND2X0_RVT U7820 ( .A1(n6700), .A2(n8161), .Y(n8405) );
  NAND2X0_RVT U7821 ( .A1(n8408), .A2(n8409), .Y(n8161) );
  NAND2X0_RVT U7822 ( .A1(n8151), .A2(n8410), .Y(n8409) );
  OR2X1_RVT U7823 ( .A1(n8150), .A2(n6706), .Y(n8410) );
  AND2X1_RVT U7824 ( .A1(n8401), .A2(n8149), .Y(n8151) );
  NAND2X0_RVT U7825 ( .A1(n6706), .A2(n8150), .Y(n8408) );
  NAND2X0_RVT U7826 ( .A1(n8411), .A2(n8412), .Y(n8150) );
  NAND2X0_RVT U7827 ( .A1(n8140), .A2(n8413), .Y(n8412) );
  OR2X1_RVT U7828 ( .A1(n8139), .A2(n6712), .Y(n8413) );
  AND2X1_RVT U7829 ( .A1(n8401), .A2(n8138), .Y(n8140) );
  NAND2X0_RVT U7830 ( .A1(n6712), .A2(n8139), .Y(n8411) );
  NAND2X0_RVT U7831 ( .A1(n8414), .A2(n8415), .Y(n8139) );
  NAND2X0_RVT U7832 ( .A1(n8129), .A2(n8416), .Y(n8415) );
  OR2X1_RVT U7833 ( .A1(n8128), .A2(n6718), .Y(n8416) );
  AND2X1_RVT U7834 ( .A1(n8401), .A2(n8417), .Y(n8129) );
  NAND2X0_RVT U7835 ( .A1(n6718), .A2(n8128), .Y(n8414) );
  NAND2X0_RVT U7836 ( .A1(n8418), .A2(n8419), .Y(n8128) );
  NAND2X0_RVT U7837 ( .A1(n8120), .A2(n8420), .Y(n8419) );
  OR2X1_RVT U7838 ( .A1(n8121), .A2(n6724), .Y(n8420) );
  AND2X1_RVT U7839 ( .A1(n8401), .A2(n8421), .Y(n8120) );
  NAND2X0_RVT U7840 ( .A1(n6739), .A2(n8422), .Y(n8401) );
  NAND2X0_RVT U7841 ( .A1(n6724), .A2(n8121), .Y(n8418) );
  NAND2X0_RVT U7842 ( .A1(n8423), .A2(n8424), .Y(n8121) );
  NAND2X0_RVT U7843 ( .A1(n8112), .A2(n6543), .Y(n8424) );
  NAND2X0_RVT U7844 ( .A1(n6543), .A2(n8107), .Y(n8423) );
  XNOR3X1_RVT U7845 ( .A1(n4931), .A2(n8112), .A3(n8425), .Y(n6543) );
  XNOR3X1_RVT U7846 ( .A1(n9575), .A2(n8426), .A3(n8427), .Y(n6724) );
  XNOR3X1_RVT U7847 ( .A1(n9569), .A2(n8428), .A3(n8429), .Y(n6718) );
  XNOR3X1_RVT U7848 ( .A1(n9566), .A2(n8430), .A3(n8431), .Y(n6712) );
  XNOR3X1_RVT U7849 ( .A1(n9565), .A2(n8432), .A3(n8433), .Y(n6706) );
  XNOR3X1_RVT U7850 ( .A1(n9564), .A2(n8434), .A3(n8435), .Y(n6700) );
  XNOR3X1_RVT U7851 ( .A1(n9563), .A2(n8436), .A3(n8437), .Y(n6694) );
  INVX0_RVT U7852 ( .A(n8185), .Y(n6688) );
  XNOR3X1_RVT U7853 ( .A1(n9562), .A2(n8192), .A3(n8438), .Y(n8185) );
  XOR2X1_RVT U7854 ( .A1(n8439), .A2(n4912), .Y(n6682) );
  XNOR2X1_RVT U7855 ( .A1(n8440), .A2(n4965), .Y(n6676) );
  NAND2X0_RVT U7856 ( .A1(n4912), .A2(n8439), .Y(n8440) );
  XNOR2X1_RVT U7857 ( .A1(n9580), .A2(n8441), .Y(n6670) );
  XNOR2X1_RVT U7858 ( .A1(n8442), .A2(n4924), .Y(n6664) );
  NAND2X0_RVT U7859 ( .A1(n8441), .A2(n4978), .Y(n8442) );
  XNOR2X1_RVT U7860 ( .A1(n9579), .A2(n8443), .Y(n6658) );
  XNOR2X1_RVT U7861 ( .A1(n8444), .A2(n4923), .Y(n6652) );
  NAND2X0_RVT U7862 ( .A1(n8443), .A2(n4977), .Y(n8444) );
  XNOR2X1_RVT U7863 ( .A1(n9578), .A2(n8445), .Y(n6646) );
  XNOR2X1_RVT U7864 ( .A1(n8446), .A2(n4922), .Y(n6640) );
  NAND2X0_RVT U7865 ( .A1(n8445), .A2(n4976), .Y(n8446) );
  XNOR2X1_RVT U7866 ( .A1(n9577), .A2(n8447), .Y(n6634) );
  XNOR2X1_RVT U7867 ( .A1(n8448), .A2(n4921), .Y(n6628) );
  NAND2X0_RVT U7868 ( .A1(n8447), .A2(n4975), .Y(n8448) );
  XNOR2X1_RVT U7869 ( .A1(n9576), .A2(n8449), .Y(n6622) );
  XNOR2X1_RVT U7870 ( .A1(n8450), .A2(n4920), .Y(n6616) );
  NAND2X0_RVT U7871 ( .A1(n8449), .A2(n4974), .Y(n8450) );
  XNOR2X1_RVT U7872 ( .A1(n9574), .A2(n8451), .Y(n6610) );
  XNOR2X1_RVT U7873 ( .A1(n8452), .A2(n4919), .Y(n6604) );
  NAND2X0_RVT U7874 ( .A1(n8451), .A2(n4973), .Y(n8452) );
  XNOR2X1_RVT U7875 ( .A1(n9573), .A2(n8453), .Y(n6598) );
  XNOR2X1_RVT U7876 ( .A1(n8454), .A2(n4918), .Y(n6592) );
  NAND2X0_RVT U7877 ( .A1(n8453), .A2(n4972), .Y(n8454) );
  XNOR2X1_RVT U7878 ( .A1(n9572), .A2(n8455), .Y(n6586) );
  XNOR2X1_RVT U7879 ( .A1(n8456), .A2(n4917), .Y(n6580) );
  NAND2X0_RVT U7880 ( .A1(n8455), .A2(n4971), .Y(n8456) );
  XNOR2X1_RVT U7881 ( .A1(n8457), .A2(n9571), .Y(n6574) );
  XNOR2X1_RVT U7882 ( .A1(n8458), .A2(n4916), .Y(n6568) );
  NAND2X0_RVT U7883 ( .A1(n8457), .A2(n4979), .Y(n8458) );
  XNOR2X1_RVT U7884 ( .A1(n8459), .A2(n9570), .Y(n6562) );
  XNOR2X1_RVT U7885 ( .A1(n8460), .A2(n4915), .Y(n6556) );
  NAND2X0_RVT U7886 ( .A1(n8459), .A2(n4970), .Y(n8460) );
  XOR2X1_RVT U7887 ( .A1(n8461), .A2(n9568), .Y(n6550) );
  XOR2X1_RVT U7888 ( .A1(n8462), .A2(n9567), .Y(n5320) );
  OR2X1_RVT U7889 ( .A1(n8461), .A2(n9568), .Y(n8462) );
  NAND3X0_RVT U7890 ( .A1(n4970), .A2(n4915), .A3(n8459), .Y(n8461) );
  AND3X1_RVT U7891 ( .A1(n4979), .A2(n4916), .A3(n8457), .Y(n8459) );
  AND3X1_RVT U7892 ( .A1(n4971), .A2(n4917), .A3(n8455), .Y(n8457) );
  AND3X1_RVT U7893 ( .A1(n4972), .A2(n4918), .A3(n8453), .Y(n8455) );
  AND3X1_RVT U7894 ( .A1(n4973), .A2(n4919), .A3(n8451), .Y(n8453) );
  AND3X1_RVT U7895 ( .A1(n4974), .A2(n4920), .A3(n8449), .Y(n8451) );
  AND3X1_RVT U7896 ( .A1(n4975), .A2(n4921), .A3(n8447), .Y(n8449) );
  AND3X1_RVT U7897 ( .A1(n4976), .A2(n4922), .A3(n8445), .Y(n8447) );
  AND3X1_RVT U7898 ( .A1(n4977), .A2(n4923), .A3(n8443), .Y(n8445) );
  AND3X1_RVT U7899 ( .A1(n4978), .A2(n4924), .A3(n8441), .Y(n8443) );
  AND3X1_RVT U7900 ( .A1(n4912), .A2(n4965), .A3(n8439), .Y(n8441) );
  NAND2X0_RVT U7901 ( .A1(n8463), .A2(n8464), .Y(n8439) );
  NAND2X0_RVT U7902 ( .A1(n8465), .A2(n5102), .Y(n8464) );
  OR2X1_RVT U7903 ( .A1(n8438), .A2(n8112), .Y(n8465) );
  NAND2X0_RVT U7904 ( .A1(n8112), .A2(n8438), .Y(n8463) );
  NAND2X0_RVT U7905 ( .A1(n8466), .A2(n8467), .Y(n8438) );
  NAND2X0_RVT U7906 ( .A1(n8468), .A2(n5103), .Y(n8467) );
  NAND2X0_RVT U7907 ( .A1(n8437), .A2(n8436), .Y(n8468) );
  OR2X1_RVT U7908 ( .A1(n8436), .A2(n8437), .Y(n8466) );
  AND2X1_RVT U7909 ( .A1(n8469), .A2(n8470), .Y(n8437) );
  NAND2X0_RVT U7910 ( .A1(n8471), .A2(n5104), .Y(n8470) );
  NAND2X0_RVT U7911 ( .A1(n8435), .A2(n8434), .Y(n8471) );
  OR2X1_RVT U7912 ( .A1(n8434), .A2(n8435), .Y(n8469) );
  AND2X1_RVT U7913 ( .A1(n8472), .A2(n8473), .Y(n8435) );
  NAND2X0_RVT U7914 ( .A1(n8474), .A2(n5105), .Y(n8473) );
  NAND2X0_RVT U7915 ( .A1(n8433), .A2(n8432), .Y(n8474) );
  OR2X1_RVT U7916 ( .A1(n8432), .A2(n8433), .Y(n8472) );
  AND2X1_RVT U7917 ( .A1(n8475), .A2(n8476), .Y(n8433) );
  NAND2X0_RVT U7918 ( .A1(n8477), .A2(n5106), .Y(n8476) );
  NAND2X0_RVT U7919 ( .A1(n8431), .A2(n8430), .Y(n8477) );
  OR2X1_RVT U7920 ( .A1(n8430), .A2(n8431), .Y(n8475) );
  AND2X1_RVT U7921 ( .A1(n8478), .A2(n8479), .Y(n8431) );
  NAND2X0_RVT U7922 ( .A1(n8480), .A2(n5107), .Y(n8479) );
  OR2X1_RVT U7923 ( .A1(n8429), .A2(n8428), .Y(n8480) );
  NAND2X0_RVT U7924 ( .A1(n8428), .A2(n8429), .Y(n8478) );
  NAND2X0_RVT U7925 ( .A1(n8481), .A2(n8482), .Y(n8429) );
  NAND2X0_RVT U7926 ( .A1(n8483), .A2(n5052), .Y(n8482) );
  OR2X1_RVT U7927 ( .A1(n8427), .A2(n8426), .Y(n8483) );
  NAND2X0_RVT U7928 ( .A1(n8426), .A2(n8427), .Y(n8481) );
  NAND2X0_RVT U7929 ( .A1(n8484), .A2(n8485), .Y(n8427) );
  NAND2X0_RVT U7930 ( .A1(n8486), .A2(n4931), .Y(n8485) );
  NAND2X0_RVT U7931 ( .A1(n8425), .A2(n8192), .Y(n8486) );
  INVX0_RVT U7932 ( .A(n8487), .Y(n8425) );
  NAND2X0_RVT U7933 ( .A1(n8112), .A2(n8487), .Y(n8484) );
  NAND4X0_RVT U7934 ( .A1(n8488), .A2(n8489), .A3(n8422), .A4(n6497), .Y(n8487) );
  NAND2X0_RVT U7935 ( .A1(n8490), .A2(n6510), .Y(n8489) );
  INVX0_RVT U7936 ( .A(n6728), .Y(n8490) );
  NAND2X0_RVT U7937 ( .A1(n8491), .A2(n6453), .Y(n6728) );
  NAND2X0_RVT U7938 ( .A1(n8112), .A2(n8107), .Y(n8488) );
  NAND4X0_RVT U7939 ( .A1(n8492), .A2(n8493), .A3(n8494), .A4(n8495), .Y(n8107) );
  NAND2X0_RVT U7940 ( .A1(n7842), .A2(n8496), .Y(n8495) );
  NAND4X0_RVT U7941 ( .A1(n8497), .A2(n8498), .A3(n8499), .A4(n8500), .Y(n8496) );
  NAND2X0_RVT U7942 ( .A1(n7694), .A2(n5123), .Y(n8500) );
  NAND2X0_RVT U7943 ( .A1(n7678), .A2(n4997), .Y(n8499) );
  NAND2X0_RVT U7944 ( .A1(n7766), .A2(n4998), .Y(n8498) );
  NAND2X0_RVT U7945 ( .A1(n8501), .A2(n4996), .Y(n8497) );
  NAND2X0_RVT U7946 ( .A1(n7853), .A2(n8502), .Y(n8494) );
  NAND2X0_RVT U7947 ( .A1(n7848), .A2(n7771), .Y(n8493) );
  NAND2X0_RVT U7948 ( .A1(n7852), .A2(n7774), .Y(n8492) );
  NAND3X0_RVT U7949 ( .A1(n8503), .A2(n8504), .A3(n6472), .Y(n8426) );
  AND2X1_RVT U7950 ( .A1(n6510), .A2(n8505), .Y(n6472) );
  NAND2X0_RVT U7951 ( .A1(n8506), .A2(n5268), .Y(n8505) );
  NAND2X0_RVT U7952 ( .A1(n8507), .A2(n8508), .Y(n8506) );
  NAND2X0_RVT U7953 ( .A1(n6739), .A2(n6742), .Y(n8508) );
  NAND2X0_RVT U7954 ( .A1(n6748), .A2(n8509), .Y(n6742) );
  NAND2X0_RVT U7955 ( .A1(n8510), .A2(n5271), .Y(n8509) );
  AND2X1_RVT U7956 ( .A1(n7010), .A2(n8511), .Y(n6748) );
  NAND4X0_RVT U7957 ( .A1(n8512), .A2(n8513), .A3(n8514), .A4(n6307), .Y(n6510) );
  NAND2X0_RVT U7958 ( .A1(n8112), .A2(n8421), .Y(n8504) );
  NAND2X0_RVT U7959 ( .A1(n6475), .A2(n8515), .Y(n8503) );
  NAND3X0_RVT U7960 ( .A1(n8422), .A2(n6497), .A3(n8516), .Y(n8428) );
  NAND2X0_RVT U7961 ( .A1(n8112), .A2(n8417), .Y(n8516) );
  NAND2X0_RVT U7962 ( .A1(n6739), .A2(n8517), .Y(n6497) );
  NAND2X0_RVT U7963 ( .A1(n8112), .A2(n8138), .Y(n8430) );
  NAND4X0_RVT U7964 ( .A1(n8518), .A2(n8519), .A3(n8520), .A4(n8521), .Y(n8138) );
  NAND2X0_RVT U7965 ( .A1(n7842), .A2(n8522), .Y(n8521) );
  NAND4X0_RVT U7966 ( .A1(n8523), .A2(n8524), .A3(n8525), .A4(n8526), .Y(n8522) );
  NAND2X0_RVT U7967 ( .A1(n7694), .A2(n5124), .Y(n8526) );
  NAND2X0_RVT U7968 ( .A1(n7678), .A2(n5017), .Y(n8525) );
  NAND2X0_RVT U7969 ( .A1(n7766), .A2(n5018), .Y(n8524) );
  NAND2X0_RVT U7970 ( .A1(n8501), .A2(n5016), .Y(n8523) );
  NAND2X0_RVT U7971 ( .A1(n7853), .A2(n8527), .Y(n8520) );
  NAND2X0_RVT U7972 ( .A1(n7848), .A2(n7719), .Y(n8519) );
  NAND2X0_RVT U7973 ( .A1(n7852), .A2(n7803), .Y(n8518) );
  NAND2X0_RVT U7974 ( .A1(n8112), .A2(n8149), .Y(n8432) );
  NAND4X0_RVT U7975 ( .A1(n8528), .A2(n8529), .A3(n8530), .A4(n8531), .Y(n8149) );
  NAND2X0_RVT U7976 ( .A1(n7842), .A2(n8532), .Y(n8531) );
  NAND4X0_RVT U7977 ( .A1(n8533), .A2(n8534), .A3(n8535), .A4(n8536), .Y(n8532) );
  NAND2X0_RVT U7978 ( .A1(n7694), .A2(n5125), .Y(n8536) );
  NAND2X0_RVT U7979 ( .A1(n7678), .A2(n5024), .Y(n8535) );
  NAND2X0_RVT U7980 ( .A1(n7766), .A2(n5025), .Y(n8534) );
  NAND2X0_RVT U7981 ( .A1(n8501), .A2(n5023), .Y(n8533) );
  NAND2X0_RVT U7982 ( .A1(n7853), .A2(n8537), .Y(n8530) );
  NAND2X0_RVT U7983 ( .A1(n7848), .A2(n7707), .Y(n8529) );
  NAND2X0_RVT U7984 ( .A1(n7852), .A2(n7813), .Y(n8528) );
  NAND2X0_RVT U7985 ( .A1(n8112), .A2(n8160), .Y(n8434) );
  NAND4X0_RVT U7986 ( .A1(n8538), .A2(n8539), .A3(n8540), .A4(n8541), .Y(n8160) );
  NAND2X0_RVT U7987 ( .A1(n7842), .A2(n8542), .Y(n8541) );
  NAND4X0_RVT U7988 ( .A1(n8543), .A2(n8544), .A3(n8545), .A4(n8546), .Y(n8542) );
  NAND2X0_RVT U7989 ( .A1(n7694), .A2(n5126), .Y(n8546) );
  NAND2X0_RVT U7990 ( .A1(n7678), .A2(n5031), .Y(n8545) );
  NAND2X0_RVT U7991 ( .A1(n7766), .A2(n5032), .Y(n8544) );
  NAND2X0_RVT U7992 ( .A1(n8501), .A2(n5030), .Y(n8543) );
  NAND2X0_RVT U7993 ( .A1(n7853), .A2(n8547), .Y(n8540) );
  NAND2X0_RVT U7994 ( .A1(n7848), .A2(n7695), .Y(n8539) );
  NAND2X0_RVT U7995 ( .A1(n7852), .A2(n7823), .Y(n8538) );
  NAND2X0_RVT U7996 ( .A1(n8112), .A2(n8171), .Y(n8436) );
  NAND4X0_RVT U7997 ( .A1(n8548), .A2(n8549), .A3(n8550), .A4(n8551), .Y(n8171) );
  NAND2X0_RVT U7998 ( .A1(n7842), .A2(n8552), .Y(n8551) );
  NAND4X0_RVT U7999 ( .A1(n8553), .A2(n8554), .A3(n8555), .A4(n8556), .Y(n8552) );
  NAND2X0_RVT U8000 ( .A1(n7694), .A2(n5127), .Y(n8556) );
  NAND2X0_RVT U8001 ( .A1(n7678), .A2(n5038), .Y(n8555) );
  NAND2X0_RVT U8002 ( .A1(n7766), .A2(n5039), .Y(n8554) );
  NAND2X0_RVT U8003 ( .A1(n8501), .A2(n5037), .Y(n8553) );
  NAND2X0_RVT U8004 ( .A1(n7853), .A2(n8557), .Y(n8550) );
  NAND2X0_RVT U8005 ( .A1(n7848), .A2(n7680), .Y(n8549) );
  NAND2X0_RVT U8006 ( .A1(n7852), .A2(n7762), .Y(n8548) );
  NAND2X0_RVT U8007 ( .A1(n8113), .A2(n5086), .Y(n8326) );
  NAND2X0_RVT U8008 ( .A1(n6731), .A2(n5380), .Y(n8558) );
  INVX0_RVT U8009 ( .A(n5479), .Y(n5380) );
  AND2X1_RVT U8010 ( .A1(n6433), .A2(n8559), .Y(n6731) );
  NAND2X0_RVT U8011 ( .A1(n5265), .A2(n6474), .Y(n8559) );
  NAND2X0_RVT U8012 ( .A1(n6434), .A2(n8422), .Y(n6474) );
  OR2X1_RVT U8013 ( .A1(n6743), .A2(n6475), .Y(n8422) );
  INVX0_RVT U8014 ( .A(n6739), .Y(n6475) );
  NAND2X0_RVT U8015 ( .A1(n7861), .A2(n5479), .Y(n8325) );
  NAND2X0_RVT U8016 ( .A1(rEIP[31]), .A2(n8114), .Y(n5315) );
  NAND4X0_RVT U8017 ( .A1(n8561), .A2(n8562), .A3(n8563), .A4(n8564), .Y(n4526) );
  NAND2X0_RVT U8018 ( .A1(n8565), .A2(n7211), .Y(n8564) );
  XNOR2X1_RVT U8019 ( .A1(n8566), .A2(n7864), .Y(n7211) );
  NAND2X0_RVT U8020 ( .A1(n8567), .A2(n4961), .Y(n8563) );
  NAND2X0_RVT U8021 ( .A1(n8568), .A2(Datao[0]), .Y(n8562) );
  NAND2X0_RVT U8022 ( .A1(n5213), .A2(n6769), .Y(n8561) );
  NAND4X0_RVT U8023 ( .A1(n8569), .A2(n8570), .A3(n8571), .A4(n8572), .Y(n4525) );
  NAND2X0_RVT U8024 ( .A1(n8565), .A2(n7231), .Y(n8572) );
  XNOR2X1_RVT U8025 ( .A1(n8573), .A2(n8574), .Y(n7231) );
  NAND2X0_RVT U8026 ( .A1(n8566), .A2(n6422), .Y(n8573) );
  NAND2X0_RVT U8027 ( .A1(n8567), .A2(n4959), .Y(n8571) );
  NAND2X0_RVT U8028 ( .A1(n8568), .A2(Datao[1]), .Y(n8570) );
  NAND2X0_RVT U8029 ( .A1(n6775), .A2(n5214), .Y(n8569) );
  NAND4X0_RVT U8030 ( .A1(n8575), .A2(n8576), .A3(n8577), .A4(n8578), .Y(n4524) );
  NAND2X0_RVT U8031 ( .A1(n8565), .A2(n7247), .Y(n8578) );
  XOR2X1_RVT U8032 ( .A1(n8579), .A2(n8580), .Y(n7247) );
  NAND2X0_RVT U8033 ( .A1(n8567), .A2(n4957), .Y(n8577) );
  NAND2X0_RVT U8034 ( .A1(n8568), .A2(Datao[2]), .Y(n8576) );
  NAND2X0_RVT U8035 ( .A1(n5212), .A2(n6781), .Y(n8575) );
  INVX0_RVT U8036 ( .A(n8581), .Y(n6781) );
  NAND4X0_RVT U8037 ( .A1(n8582), .A2(n8583), .A3(n8584), .A4(n8585), .Y(n4523) );
  NAND2X0_RVT U8038 ( .A1(n8565), .A2(n7280), .Y(n8585) );
  XNOR2X1_RVT U8039 ( .A1(n8586), .A2(n8587), .Y(n7280) );
  NAND2X0_RVT U8040 ( .A1(n8579), .A2(n8580), .Y(n8586) );
  NAND2X0_RVT U8041 ( .A1(n8567), .A2(n4951), .Y(n8584) );
  NAND2X0_RVT U8042 ( .A1(n8568), .A2(Datao[3]), .Y(n8583) );
  NAND2X0_RVT U8043 ( .A1(n5215), .A2(n6787), .Y(n8582) );
  INVX0_RVT U8044 ( .A(n8588), .Y(n6787) );
  NAND4X0_RVT U8045 ( .A1(n8589), .A2(n8590), .A3(n8591), .A4(n8592), .Y(n4522) );
  NAND2X0_RVT U8046 ( .A1(n8565), .A2(n7291), .Y(n8592) );
  XOR2X1_RVT U8047 ( .A1(n8593), .A2(n8594), .Y(n7291) );
  NAND2X0_RVT U8048 ( .A1(n8567), .A2(n4954), .Y(n8591) );
  NAND2X0_RVT U8049 ( .A1(n8568), .A2(Datao[4]), .Y(n8590) );
  NAND2X0_RVT U8050 ( .A1(n5214), .A2(n6793), .Y(n8589) );
  INVX0_RVT U8051 ( .A(n8595), .Y(n6793) );
  NAND4X0_RVT U8052 ( .A1(n8596), .A2(n8597), .A3(n8598), .A4(n8599), .Y(n4521) );
  NAND2X0_RVT U8053 ( .A1(n8565), .A2(n7302), .Y(n8599) );
  XNOR2X1_RVT U8054 ( .A1(n8600), .A2(n8601), .Y(n7302) );
  NAND2X0_RVT U8055 ( .A1(n8593), .A2(n8594), .Y(n8600) );
  NAND2X0_RVT U8056 ( .A1(n8567), .A2(n4948), .Y(n8598) );
  NAND2X0_RVT U8057 ( .A1(n8568), .A2(Datao[5]), .Y(n8597) );
  NAND2X0_RVT U8058 ( .A1(n5213), .A2(n6799), .Y(n8596) );
  INVX0_RVT U8059 ( .A(n8602), .Y(n6799) );
  NAND4X0_RVT U8060 ( .A1(n8603), .A2(n8604), .A3(n8605), .A4(n8606), .Y(n4520) );
  NAND2X0_RVT U8061 ( .A1(n8565), .A2(n7313), .Y(n8606) );
  XOR2X1_RVT U8062 ( .A1(n8607), .A2(n8608), .Y(n7313) );
  NAND2X0_RVT U8063 ( .A1(n8567), .A2(n4956), .Y(n8605) );
  NAND2X0_RVT U8064 ( .A1(n8568), .A2(Datao[6]), .Y(n8604) );
  NAND2X0_RVT U8065 ( .A1(n5212), .A2(n6805), .Y(n8603) );
  INVX0_RVT U8066 ( .A(n8609), .Y(n6805) );
  NAND4X0_RVT U8067 ( .A1(n8610), .A2(n8611), .A3(n8612), .A4(n8613), .Y(n4519) );
  NAND2X0_RVT U8068 ( .A1(n8565), .A2(n7324), .Y(n8613) );
  XNOR2X1_RVT U8069 ( .A1(n8614), .A2(n8615), .Y(n7324) );
  NAND2X0_RVT U8070 ( .A1(n8607), .A2(n8608), .Y(n8614) );
  NAND2X0_RVT U8071 ( .A1(n8567), .A2(n4950), .Y(n8612) );
  NAND2X0_RVT U8072 ( .A1(n8568), .A2(Datao[7]), .Y(n8611) );
  NAND2X0_RVT U8073 ( .A1(n5215), .A2(n6811), .Y(n8610) );
  INVX0_RVT U8074 ( .A(n8616), .Y(n6811) );
  NAND4X0_RVT U8075 ( .A1(n8617), .A2(n8618), .A3(n8619), .A4(n8620), .Y(n4518) );
  NAND2X0_RVT U8076 ( .A1(n8565), .A2(n7335), .Y(n8620) );
  XOR2X1_RVT U8077 ( .A1(n8621), .A2(n8622), .Y(n7335) );
  NAND2X0_RVT U8078 ( .A1(n8567), .A2(n4953), .Y(n8619) );
  NAND2X0_RVT U8079 ( .A1(n8568), .A2(Datao[8]), .Y(n8618) );
  NAND2X0_RVT U8080 ( .A1(n5214), .A2(n6817), .Y(n8617) );
  INVX0_RVT U8081 ( .A(n8623), .Y(n6817) );
  NAND4X0_RVT U8082 ( .A1(n8624), .A2(n8625), .A3(n8626), .A4(n8627), .Y(n4517) );
  NAND2X0_RVT U8083 ( .A1(n8565), .A2(n7346), .Y(n8627) );
  XNOR2X1_RVT U8084 ( .A1(n8628), .A2(n8629), .Y(n7346) );
  NAND2X0_RVT U8085 ( .A1(n8621), .A2(n8622), .Y(n8628) );
  NAND2X0_RVT U8086 ( .A1(n8567), .A2(n4947), .Y(n8626) );
  NAND2X0_RVT U8087 ( .A1(n8568), .A2(Datao[9]), .Y(n8625) );
  NAND2X0_RVT U8088 ( .A1(n5213), .A2(n6823), .Y(n8624) );
  INVX0_RVT U8089 ( .A(n8630), .Y(n6823) );
  NAND4X0_RVT U8090 ( .A1(n8631), .A2(n8632), .A3(n8633), .A4(n8634), .Y(n4516) );
  NAND2X0_RVT U8091 ( .A1(n8565), .A2(n7357), .Y(n8634) );
  XOR2X1_RVT U8092 ( .A1(n8635), .A2(n8636), .Y(n7357) );
  NAND2X0_RVT U8093 ( .A1(n8567), .A2(n4952), .Y(n8633) );
  NAND2X0_RVT U8094 ( .A1(n8568), .A2(Datao[10]), .Y(n8632) );
  NAND2X0_RVT U8095 ( .A1(n5212), .A2(n6829), .Y(n8631) );
  INVX0_RVT U8096 ( .A(n8637), .Y(n6829) );
  NAND4X0_RVT U8097 ( .A1(n8638), .A2(n8639), .A3(n8640), .A4(n8641), .Y(n4515) );
  NAND2X0_RVT U8098 ( .A1(n8565), .A2(n7368), .Y(n8641) );
  XNOR2X1_RVT U8099 ( .A1(n8642), .A2(n8643), .Y(n7368) );
  NAND2X0_RVT U8100 ( .A1(n8635), .A2(n8636), .Y(n8642) );
  NAND2X0_RVT U8101 ( .A1(n8567), .A2(n4946), .Y(n8640) );
  NAND2X0_RVT U8102 ( .A1(n8568), .A2(Datao[11]), .Y(n8639) );
  NAND2X0_RVT U8103 ( .A1(n5215), .A2(n6835), .Y(n8638) );
  INVX0_RVT U8104 ( .A(n8644), .Y(n6835) );
  NAND4X0_RVT U8105 ( .A1(n8645), .A2(n8646), .A3(n8647), .A4(n8648), .Y(n4514) );
  NAND2X0_RVT U8106 ( .A1(n8565), .A2(n7379), .Y(n8648) );
  XOR2X1_RVT U8107 ( .A1(n8649), .A2(n8650), .Y(n7379) );
  NAND2X0_RVT U8108 ( .A1(n8567), .A2(n4955), .Y(n8647) );
  NAND2X0_RVT U8109 ( .A1(n8568), .A2(Datao[12]), .Y(n8646) );
  NAND2X0_RVT U8110 ( .A1(n5214), .A2(n6841), .Y(n8645) );
  INVX0_RVT U8111 ( .A(n8651), .Y(n6841) );
  NAND4X0_RVT U8112 ( .A1(n8652), .A2(n8653), .A3(n8654), .A4(n8655), .Y(n4513) );
  NAND2X0_RVT U8113 ( .A1(n8565), .A2(n7390), .Y(n8655) );
  XNOR2X1_RVT U8114 ( .A1(n8656), .A2(n8657), .Y(n7390) );
  NAND2X0_RVT U8115 ( .A1(n8649), .A2(n8650), .Y(n8656) );
  NAND2X0_RVT U8116 ( .A1(n8567), .A2(n4949), .Y(n8654) );
  NAND2X0_RVT U8117 ( .A1(n8568), .A2(Datao[13]), .Y(n8653) );
  NAND2X0_RVT U8118 ( .A1(n5213), .A2(n6847), .Y(n8652) );
  INVX0_RVT U8119 ( .A(n8658), .Y(n6847) );
  NAND4X0_RVT U8120 ( .A1(n8659), .A2(n8660), .A3(n8661), .A4(n8662), .Y(n4512) );
  NAND2X0_RVT U8121 ( .A1(n8565), .A2(n7401), .Y(n8662) );
  XOR2X1_RVT U8122 ( .A1(n8663), .A2(n8664), .Y(n7401) );
  NAND2X0_RVT U8123 ( .A1(n8567), .A2(n4960), .Y(n8661) );
  NAND2X0_RVT U8124 ( .A1(n8568), .A2(Datao[14]), .Y(n8660) );
  NAND2X0_RVT U8125 ( .A1(n5212), .A2(n6853), .Y(n8659) );
  NAND4X0_RVT U8126 ( .A1(n8665), .A2(n8666), .A3(n8667), .A4(n8668), .Y(n4511) );
  NAND2X0_RVT U8127 ( .A1(n5215), .A2(n6859), .Y(n8668) );
  NAND2X0_RVT U8128 ( .A1(n8669), .A2(n8670), .Y(n6859) );
  NAND2X0_RVT U8129 ( .A1(n5214), .A2(n5174), .Y(n8670) );
  XNOR2X1_RVT U8130 ( .A1(n8671), .A2(n8672), .Y(n8669) );
  NAND2X0_RVT U8131 ( .A1(n8567), .A2(n4945), .Y(n8667) );
  AND3X1_RVT U8132 ( .A1(n5265), .A2(n8673), .A3(n8510), .Y(n8567) );
  NAND2X0_RVT U8133 ( .A1(n8565), .A2(n7412), .Y(n8666) );
  XOR2X1_RVT U8134 ( .A1(n8674), .A2(n8675), .Y(n7412) );
  NAND2X0_RVT U8135 ( .A1(n8568), .A2(Datao[15]), .Y(n8665) );
  NAND3X0_RVT U8136 ( .A1(n8676), .A2(n8677), .A3(n8678), .Y(n4510) );
  NAND2X0_RVT U8137 ( .A1(n8568), .A2(Datao[16]), .Y(n8678) );
  NAND2X0_RVT U8138 ( .A1(n5213), .A2(n6916), .Y(n8677) );
  XOR2X1_RVT U8139 ( .A1(n8679), .A2(n8680), .Y(n6916) );
  NAND2X0_RVT U8140 ( .A1(n8565), .A2(n7423), .Y(n8676) );
  XOR2X1_RVT U8141 ( .A1(n8681), .A2(n8682), .Y(n7423) );
  OR2X1_RVT U8142 ( .A1(n6769), .A2(n8683), .Y(n8681) );
  XOR2X1_RVT U8143 ( .A1(n8684), .A2(n8685), .Y(n6769) );
  NAND3X0_RVT U8144 ( .A1(n8686), .A2(n8687), .A3(n8688), .Y(n4509) );
  NAND2X0_RVT U8145 ( .A1(n8568), .A2(Datao[17]), .Y(n8688) );
  NAND2X0_RVT U8146 ( .A1(n5212), .A2(n6922), .Y(n8687) );
  XOR2X1_RVT U8147 ( .A1(n8689), .A2(n8690), .Y(n6922) );
  NAND2X0_RVT U8148 ( .A1(n8565), .A2(n7440), .Y(n8686) );
  XOR2X1_RVT U8149 ( .A1(n8691), .A2(n8692), .Y(n7440) );
  OR2X1_RVT U8150 ( .A1(n6775), .A2(n8693), .Y(n8691) );
  XNOR3X1_RVT U8151 ( .A1(n8694), .A2(n8695), .A3(n8696), .Y(n6775) );
  NAND3X0_RVT U8152 ( .A1(n8697), .A2(n8698), .A3(n8699), .Y(n4508) );
  NAND2X0_RVT U8153 ( .A1(n8568), .A2(Datao[18]), .Y(n8699) );
  NAND2X0_RVT U8154 ( .A1(n5215), .A2(n6928), .Y(n8698) );
  XOR2X1_RVT U8155 ( .A1(n8700), .A2(n8701), .Y(n6928) );
  NAND2X0_RVT U8156 ( .A1(n8565), .A2(n7456), .Y(n8697) );
  XOR2X1_RVT U8157 ( .A1(n8702), .A2(n8703), .Y(n7456) );
  NAND2X0_RVT U8158 ( .A1(n8581), .A2(n8704), .Y(n8702) );
  XNOR3X1_RVT U8159 ( .A1(n8705), .A2(n8706), .A3(n8707), .Y(n8581) );
  NAND3X0_RVT U8160 ( .A1(n8708), .A2(n8709), .A3(n8710), .Y(n4507) );
  NAND2X0_RVT U8161 ( .A1(n8568), .A2(Datao[19]), .Y(n8710) );
  NAND2X0_RVT U8162 ( .A1(n5214), .A2(n6934), .Y(n8709) );
  XOR2X1_RVT U8163 ( .A1(n8711), .A2(n8712), .Y(n6934) );
  NAND2X0_RVT U8164 ( .A1(n8565), .A2(n7472), .Y(n8708) );
  XOR2X1_RVT U8165 ( .A1(n8713), .A2(n8714), .Y(n7472) );
  NAND2X0_RVT U8166 ( .A1(n8588), .A2(n8715), .Y(n8713) );
  XNOR3X1_RVT U8167 ( .A1(n8716), .A2(n8717), .A3(n8718), .Y(n8588) );
  NAND3X0_RVT U8168 ( .A1(n8719), .A2(n8720), .A3(n8721), .Y(n4506) );
  NAND2X0_RVT U8169 ( .A1(n8568), .A2(Datao[20]), .Y(n8721) );
  NAND2X0_RVT U8170 ( .A1(n5213), .A2(n6940), .Y(n8720) );
  XOR2X1_RVT U8171 ( .A1(n8722), .A2(n8723), .Y(n6940) );
  NAND2X0_RVT U8172 ( .A1(n8565), .A2(n7489), .Y(n8719) );
  XOR2X1_RVT U8173 ( .A1(n8724), .A2(n8725), .Y(n7489) );
  NAND2X0_RVT U8174 ( .A1(n8595), .A2(n8726), .Y(n8724) );
  XNOR3X1_RVT U8175 ( .A1(n8727), .A2(n8728), .A3(n8729), .Y(n8595) );
  NAND3X0_RVT U8176 ( .A1(n8730), .A2(n8731), .A3(n8732), .Y(n4505) );
  NAND2X0_RVT U8177 ( .A1(n8568), .A2(Datao[21]), .Y(n8732) );
  NAND2X0_RVT U8178 ( .A1(n5212), .A2(n6946), .Y(n8731) );
  XOR2X1_RVT U8179 ( .A1(n8733), .A2(n8734), .Y(n6946) );
  NAND2X0_RVT U8180 ( .A1(n8565), .A2(n7505), .Y(n8730) );
  XOR2X1_RVT U8181 ( .A1(n8735), .A2(n8736), .Y(n7505) );
  NAND2X0_RVT U8182 ( .A1(n8602), .A2(n8737), .Y(n8735) );
  XNOR3X1_RVT U8183 ( .A1(n8738), .A2(n8739), .A3(n8740), .Y(n8602) );
  NAND3X0_RVT U8184 ( .A1(n8741), .A2(n8742), .A3(n8743), .Y(n4504) );
  NAND2X0_RVT U8185 ( .A1(n8568), .A2(Datao[22]), .Y(n8743) );
  NAND2X0_RVT U8186 ( .A1(n5215), .A2(n6952), .Y(n8742) );
  XOR2X1_RVT U8187 ( .A1(n8744), .A2(n8745), .Y(n6952) );
  NAND2X0_RVT U8188 ( .A1(n8565), .A2(n7521), .Y(n8741) );
  XOR2X1_RVT U8189 ( .A1(n8746), .A2(n8747), .Y(n7521) );
  NAND2X0_RVT U8190 ( .A1(n8609), .A2(n8748), .Y(n8746) );
  XNOR3X1_RVT U8191 ( .A1(n8749), .A2(n8750), .A3(n8751), .Y(n8609) );
  NAND3X0_RVT U8192 ( .A1(n8752), .A2(n8753), .A3(n8754), .Y(n4503) );
  NAND2X0_RVT U8193 ( .A1(n8568), .A2(Datao[23]), .Y(n8754) );
  NAND2X0_RVT U8194 ( .A1(n5214), .A2(n6958), .Y(n8753) );
  XOR2X1_RVT U8195 ( .A1(n8755), .A2(n8756), .Y(n6958) );
  NAND2X0_RVT U8196 ( .A1(n8565), .A2(n7537), .Y(n8752) );
  XOR2X1_RVT U8197 ( .A1(n8757), .A2(n8758), .Y(n7537) );
  NAND2X0_RVT U8198 ( .A1(n8616), .A2(n8759), .Y(n8757) );
  XNOR3X1_RVT U8199 ( .A1(n8760), .A2(n8761), .A3(n8762), .Y(n8616) );
  NAND3X0_RVT U8200 ( .A1(n8763), .A2(n8764), .A3(n8765), .Y(n4502) );
  NAND2X0_RVT U8201 ( .A1(n8568), .A2(Datao[24]), .Y(n8765) );
  NAND2X0_RVT U8202 ( .A1(n5213), .A2(n6964), .Y(n8764) );
  XOR2X1_RVT U8203 ( .A1(n8766), .A2(n8767), .Y(n6964) );
  NAND2X0_RVT U8204 ( .A1(n8565), .A2(n7554), .Y(n8763) );
  XOR2X1_RVT U8205 ( .A1(n8768), .A2(n8769), .Y(n7554) );
  NAND2X0_RVT U8206 ( .A1(n8623), .A2(n8770), .Y(n8768) );
  XNOR3X1_RVT U8207 ( .A1(n8771), .A2(n8772), .A3(n8773), .Y(n8623) );
  NAND3X0_RVT U8208 ( .A1(n8774), .A2(n8775), .A3(n8776), .Y(n4501) );
  NAND2X0_RVT U8209 ( .A1(n8568), .A2(Datao[25]), .Y(n8776) );
  NAND2X0_RVT U8210 ( .A1(n5212), .A2(n6970), .Y(n8775) );
  XOR2X1_RVT U8211 ( .A1(n8777), .A2(n8778), .Y(n6970) );
  NAND2X0_RVT U8212 ( .A1(n8565), .A2(n7572), .Y(n8774) );
  XOR2X1_RVT U8213 ( .A1(n8779), .A2(n8780), .Y(n7572) );
  NAND2X0_RVT U8214 ( .A1(n8630), .A2(n8781), .Y(n8779) );
  XNOR3X1_RVT U8215 ( .A1(n8782), .A2(n8783), .A3(n8784), .Y(n8630) );
  NAND3X0_RVT U8216 ( .A1(n8785), .A2(n8786), .A3(n8787), .Y(n4500) );
  NAND2X0_RVT U8217 ( .A1(n8568), .A2(Datao[26]), .Y(n8787) );
  NAND2X0_RVT U8218 ( .A1(n5215), .A2(n6976), .Y(n8786) );
  XOR2X1_RVT U8219 ( .A1(n8788), .A2(n8789), .Y(n6976) );
  NAND2X0_RVT U8220 ( .A1(n8565), .A2(n7590), .Y(n8785) );
  XOR2X1_RVT U8221 ( .A1(n8790), .A2(n8791), .Y(n7590) );
  NAND2X0_RVT U8222 ( .A1(n8637), .A2(n8792), .Y(n8790) );
  XNOR3X1_RVT U8223 ( .A1(n8793), .A2(n8794), .A3(n8795), .Y(n8637) );
  NAND3X0_RVT U8224 ( .A1(n8796), .A2(n8797), .A3(n8798), .Y(n4499) );
  NAND2X0_RVT U8225 ( .A1(n8568), .A2(Datao[27]), .Y(n8798) );
  NAND2X0_RVT U8226 ( .A1(n5214), .A2(n6982), .Y(n8797) );
  XOR2X1_RVT U8227 ( .A1(n8799), .A2(n8800), .Y(n6982) );
  NAND2X0_RVT U8228 ( .A1(n8565), .A2(n7608), .Y(n8796) );
  XOR2X1_RVT U8229 ( .A1(n8801), .A2(n8802), .Y(n7608) );
  NAND2X0_RVT U8230 ( .A1(n8644), .A2(n8803), .Y(n8801) );
  XNOR3X1_RVT U8231 ( .A1(n8804), .A2(n8805), .A3(n8806), .Y(n8644) );
  NAND3X0_RVT U8232 ( .A1(n8807), .A2(n8808), .A3(n8809), .Y(n4498) );
  NAND2X0_RVT U8233 ( .A1(n8568), .A2(Datao[28]), .Y(n8809) );
  NAND2X0_RVT U8234 ( .A1(n5213), .A2(n6988), .Y(n8808) );
  XOR2X1_RVT U8235 ( .A1(n8810), .A2(n8811), .Y(n6988) );
  NAND2X0_RVT U8236 ( .A1(n8565), .A2(n7626), .Y(n8807) );
  XOR2X1_RVT U8237 ( .A1(n8812), .A2(n8813), .Y(n7626) );
  NAND2X0_RVT U8238 ( .A1(n8651), .A2(n8814), .Y(n8812) );
  XNOR3X1_RVT U8239 ( .A1(n8815), .A2(n8816), .A3(n8817), .Y(n8651) );
  NAND3X0_RVT U8240 ( .A1(n8818), .A2(n8819), .A3(n8820), .Y(n4497) );
  NAND2X0_RVT U8241 ( .A1(n8568), .A2(Datao[29]), .Y(n8820) );
  NAND2X0_RVT U8242 ( .A1(n5212), .A2(n6994), .Y(n8819) );
  XOR2X1_RVT U8243 ( .A1(n8821), .A2(n8822), .Y(n6994) );
  NAND2X0_RVT U8244 ( .A1(n8565), .A2(n7644), .Y(n8818) );
  XOR2X1_RVT U8245 ( .A1(n8823), .A2(n8824), .Y(n7644) );
  NAND2X0_RVT U8246 ( .A1(n8658), .A2(n8825), .Y(n8823) );
  XNOR3X1_RVT U8247 ( .A1(n8826), .A2(n8827), .A3(n8828), .Y(n8658) );
  NAND3X0_RVT U8248 ( .A1(n8829), .A2(n8830), .A3(n8831), .Y(n4496) );
  NAND2X0_RVT U8249 ( .A1(n8568), .A2(Datao[30]), .Y(n8831) );
  NAND2X0_RVT U8250 ( .A1(n5215), .A2(n7000), .Y(n8830) );
  XOR2X1_RVT U8251 ( .A1(n7013), .A2(n7014), .Y(n7000) );
  NAND2X0_RVT U8252 ( .A1(n8832), .A2(n8833), .Y(n7014) );
  NAND2X0_RVT U8253 ( .A1(n5206), .A2(n5101), .Y(n8833) );
  NAND2X0_RVT U8254 ( .A1(uWord[14]), .A2(n5213), .Y(n8832) );
  AND2X1_RVT U8255 ( .A1(n8821), .A2(n8822), .Y(n7013) );
  NAND2X0_RVT U8256 ( .A1(n8834), .A2(n8835), .Y(n8822) );
  NAND2X0_RVT U8257 ( .A1(n5205), .A2(n5100), .Y(n8835) );
  NAND2X0_RVT U8258 ( .A1(uWord[13]), .A2(n5212), .Y(n8834) );
  AND2X1_RVT U8259 ( .A1(n8810), .A2(n8811), .Y(n8821) );
  NAND2X0_RVT U8260 ( .A1(n8836), .A2(n8837), .Y(n8811) );
  NAND2X0_RVT U8261 ( .A1(n5204), .A2(n5099), .Y(n8837) );
  NAND2X0_RVT U8262 ( .A1(uWord[12]), .A2(n5215), .Y(n8836) );
  AND2X1_RVT U8263 ( .A1(n8799), .A2(n8800), .Y(n8810) );
  NAND2X0_RVT U8264 ( .A1(n8838), .A2(n8839), .Y(n8800) );
  NAND2X0_RVT U8265 ( .A1(n5207), .A2(n5098), .Y(n8839) );
  NAND2X0_RVT U8266 ( .A1(uWord[11]), .A2(n5214), .Y(n8838) );
  AND2X1_RVT U8267 ( .A1(n8788), .A2(n8789), .Y(n8799) );
  NAND2X0_RVT U8268 ( .A1(n8840), .A2(n8841), .Y(n8789) );
  NAND2X0_RVT U8269 ( .A1(n5206), .A2(n5097), .Y(n8841) );
  NAND2X0_RVT U8270 ( .A1(uWord[10]), .A2(n5213), .Y(n8840) );
  AND2X1_RVT U8271 ( .A1(n8777), .A2(n8778), .Y(n8788) );
  NAND2X0_RVT U8272 ( .A1(n8842), .A2(n8843), .Y(n8778) );
  NAND2X0_RVT U8273 ( .A1(n5205), .A2(n5096), .Y(n8843) );
  NAND2X0_RVT U8274 ( .A1(uWord[9]), .A2(n5212), .Y(n8842) );
  AND2X1_RVT U8275 ( .A1(n8766), .A2(n8767), .Y(n8777) );
  NAND2X0_RVT U8276 ( .A1(n8844), .A2(n8845), .Y(n8767) );
  NAND2X0_RVT U8277 ( .A1(n5204), .A2(n5095), .Y(n8845) );
  NAND2X0_RVT U8278 ( .A1(uWord[8]), .A2(n5215), .Y(n8844) );
  AND2X1_RVT U8279 ( .A1(n8755), .A2(n8756), .Y(n8766) );
  NAND2X0_RVT U8280 ( .A1(n8846), .A2(n8847), .Y(n8756) );
  NAND2X0_RVT U8281 ( .A1(n5207), .A2(n5094), .Y(n8847) );
  NAND2X0_RVT U8282 ( .A1(uWord[7]), .A2(n5214), .Y(n8846) );
  AND2X1_RVT U8283 ( .A1(n8744), .A2(n8745), .Y(n8755) );
  NAND2X0_RVT U8284 ( .A1(n8848), .A2(n8849), .Y(n8745) );
  NAND2X0_RVT U8285 ( .A1(n5206), .A2(n5093), .Y(n8849) );
  NAND2X0_RVT U8286 ( .A1(uWord[6]), .A2(n5213), .Y(n8848) );
  AND2X1_RVT U8287 ( .A1(n8733), .A2(n8734), .Y(n8744) );
  NAND2X0_RVT U8288 ( .A1(n8850), .A2(n8851), .Y(n8734) );
  NAND2X0_RVT U8289 ( .A1(n5205), .A2(n5092), .Y(n8851) );
  NAND2X0_RVT U8290 ( .A1(uWord[5]), .A2(n5212), .Y(n8850) );
  AND2X1_RVT U8291 ( .A1(n8722), .A2(n8723), .Y(n8733) );
  NAND2X0_RVT U8292 ( .A1(n8852), .A2(n8853), .Y(n8723) );
  NAND2X0_RVT U8293 ( .A1(n5204), .A2(n5091), .Y(n8853) );
  NAND2X0_RVT U8294 ( .A1(uWord[4]), .A2(n5215), .Y(n8852) );
  AND2X1_RVT U8295 ( .A1(n8711), .A2(n8712), .Y(n8722) );
  NAND2X0_RVT U8296 ( .A1(n8854), .A2(n8855), .Y(n8712) );
  NAND2X0_RVT U8297 ( .A1(n5207), .A2(n5090), .Y(n8855) );
  NAND2X0_RVT U8298 ( .A1(uWord[3]), .A2(n5214), .Y(n8854) );
  AND2X1_RVT U8299 ( .A1(n8700), .A2(n8701), .Y(n8711) );
  NAND2X0_RVT U8300 ( .A1(n8856), .A2(n8857), .Y(n8701) );
  NAND2X0_RVT U8301 ( .A1(n5206), .A2(n5089), .Y(n8857) );
  NAND2X0_RVT U8302 ( .A1(uWord[2]), .A2(n5213), .Y(n8856) );
  AND2X1_RVT U8303 ( .A1(n8689), .A2(n8690), .Y(n8700) );
  NAND2X0_RVT U8304 ( .A1(n8858), .A2(n8859), .Y(n8690) );
  NAND2X0_RVT U8305 ( .A1(n5205), .A2(n5087), .Y(n8859) );
  NAND2X0_RVT U8306 ( .A1(uWord[1]), .A2(n5212), .Y(n8858) );
  AND2X1_RVT U8307 ( .A1(n8679), .A2(n8680), .Y(n8689) );
  NAND2X0_RVT U8308 ( .A1(n8860), .A2(n8861), .Y(n8680) );
  NAND2X0_RVT U8309 ( .A1(n5204), .A2(n5088), .Y(n8861) );
  NAND2X0_RVT U8310 ( .A1(uWord[0]), .A2(n5215), .Y(n8860) );
  AND2X1_RVT U8311 ( .A1(n8672), .A2(n8671), .Y(n8679) );
  AND2X1_RVT U8312 ( .A1(n8862), .A2(n8863), .Y(n8671) );
  INVX0_RVT U8313 ( .A(n8864), .Y(n8862) );
  AND2X1_RVT U8314 ( .A1(n5204), .A2(n4945), .Y(n8672) );
  NAND2X0_RVT U8315 ( .A1(n8565), .A2(n7662), .Y(n8829) );
  XOR2X1_RVT U8316 ( .A1(n8865), .A2(n7909), .Y(n7662) );
  AND2X1_RVT U8317 ( .A1(n8866), .A2(n8824), .Y(n7909) );
  AND2X1_RVT U8318 ( .A1(n8867), .A2(n8813), .Y(n8824) );
  AND2X1_RVT U8319 ( .A1(n8868), .A2(n8802), .Y(n8813) );
  AND2X1_RVT U8320 ( .A1(n8869), .A2(n8791), .Y(n8802) );
  AND2X1_RVT U8321 ( .A1(n8870), .A2(n8780), .Y(n8791) );
  AND2X1_RVT U8322 ( .A1(n8871), .A2(n8769), .Y(n8780) );
  AND2X1_RVT U8323 ( .A1(n8872), .A2(n8758), .Y(n8769) );
  AND2X1_RVT U8324 ( .A1(n8873), .A2(n8747), .Y(n8758) );
  AND2X1_RVT U8325 ( .A1(n8874), .A2(n8736), .Y(n8747) );
  AND2X1_RVT U8326 ( .A1(n8875), .A2(n8725), .Y(n8736) );
  AND2X1_RVT U8327 ( .A1(n8876), .A2(n8714), .Y(n8725) );
  AND2X1_RVT U8328 ( .A1(n8877), .A2(n8703), .Y(n8714) );
  AND2X1_RVT U8329 ( .A1(n8693), .A2(n8692), .Y(n8703) );
  AND2X1_RVT U8330 ( .A1(n8683), .A2(n8682), .Y(n8692) );
  AND2X1_RVT U8331 ( .A1(n9537), .A2(n6422), .Y(n8682) );
  AND2X1_RVT U8332 ( .A1(n8674), .A2(n8675), .Y(n8683) );
  XNOR2X1_RVT U8333 ( .A1(n8878), .A2(n7864), .Y(n8675) );
  NAND2X0_RVT U8334 ( .A1(n8879), .A2(n8880), .Y(n8878) );
  NAND2X0_RVT U8335 ( .A1(n6422), .A2(n4932), .Y(n8880) );
  NAND2X0_RVT U8336 ( .A1(n8881), .A2(n4945), .Y(n8879) );
  AND2X1_RVT U8337 ( .A1(n8663), .A2(n8664), .Y(n8674) );
  XNOR2X1_RVT U8338 ( .A1(n8882), .A2(n7864), .Y(n8664) );
  NAND2X0_RVT U8339 ( .A1(n8883), .A2(n8884), .Y(n8882) );
  NAND2X0_RVT U8340 ( .A1(n6422), .A2(n4934), .Y(n8884) );
  NAND2X0_RVT U8341 ( .A1(n8881), .A2(n4960), .Y(n8883) );
  AND3X1_RVT U8342 ( .A1(n8650), .A2(n8649), .A3(n8657), .Y(n8663) );
  XNOR2X1_RVT U8343 ( .A1(n8885), .A2(n7864), .Y(n8657) );
  NAND2X0_RVT U8344 ( .A1(n8886), .A2(n8887), .Y(n8885) );
  NAND2X0_RVT U8345 ( .A1(n6422), .A2(n4935), .Y(n8887) );
  NAND2X0_RVT U8346 ( .A1(n8881), .A2(n4949), .Y(n8886) );
  AND3X1_RVT U8347 ( .A1(n8636), .A2(n8635), .A3(n8643), .Y(n8649) );
  XNOR2X1_RVT U8348 ( .A1(n8888), .A2(n7864), .Y(n8643) );
  NAND2X0_RVT U8349 ( .A1(n8889), .A2(n8890), .Y(n8888) );
  NAND2X0_RVT U8350 ( .A1(n6422), .A2(n4936), .Y(n8890) );
  NAND2X0_RVT U8351 ( .A1(n8881), .A2(n4946), .Y(n8889) );
  AND3X1_RVT U8352 ( .A1(n8622), .A2(n8621), .A3(n8629), .Y(n8635) );
  XNOR2X1_RVT U8353 ( .A1(n8891), .A2(n7864), .Y(n8629) );
  NAND2X0_RVT U8354 ( .A1(n8892), .A2(n8893), .Y(n8891) );
  NAND2X0_RVT U8355 ( .A1(n6422), .A2(n4933), .Y(n8893) );
  NAND2X0_RVT U8356 ( .A1(n8881), .A2(n4947), .Y(n8892) );
  AND3X1_RVT U8357 ( .A1(n8608), .A2(n8607), .A3(n8615), .Y(n8621) );
  XNOR2X1_RVT U8358 ( .A1(n8894), .A2(n7864), .Y(n8615) );
  NAND2X0_RVT U8359 ( .A1(n8895), .A2(n8896), .Y(n8894) );
  NAND2X0_RVT U8360 ( .A1(n6422), .A2(n4937), .Y(n8896) );
  NAND2X0_RVT U8361 ( .A1(n8881), .A2(n4950), .Y(n8895) );
  AND3X1_RVT U8362 ( .A1(n8594), .A2(n8593), .A3(n8601), .Y(n8607) );
  XNOR2X1_RVT U8363 ( .A1(n8897), .A2(n7864), .Y(n8601) );
  NAND2X0_RVT U8364 ( .A1(n8898), .A2(n8899), .Y(n8897) );
  NAND2X0_RVT U8365 ( .A1(n6422), .A2(n4938), .Y(n8899) );
  NAND2X0_RVT U8366 ( .A1(n8881), .A2(n4948), .Y(n8898) );
  AND3X1_RVT U8367 ( .A1(n8580), .A2(n8579), .A3(n8587), .Y(n8593) );
  XNOR2X1_RVT U8368 ( .A1(n8900), .A2(n7864), .Y(n8587) );
  NAND2X0_RVT U8369 ( .A1(n8901), .A2(n8902), .Y(n8900) );
  NAND2X0_RVT U8370 ( .A1(n6422), .A2(n4939), .Y(n8902) );
  NAND2X0_RVT U8371 ( .A1(n8881), .A2(n4951), .Y(n8901) );
  AND3X1_RVT U8372 ( .A1(n8566), .A2(n6422), .A3(n8574), .Y(n8579) );
  XNOR2X1_RVT U8373 ( .A1(n8903), .A2(n7864), .Y(n8574) );
  NAND2X0_RVT U8374 ( .A1(n8904), .A2(n8905), .Y(n8903) );
  NAND2X0_RVT U8375 ( .A1(n6422), .A2(n4964), .Y(n8905) );
  NAND2X0_RVT U8376 ( .A1(n8881), .A2(n4959), .Y(n8904) );
  XOR2X1_RVT U8377 ( .A1(n8906), .A2(n6422), .Y(n8566) );
  NAND2X0_RVT U8378 ( .A1(n8907), .A2(n8908), .Y(n8906) );
  NAND2X0_RVT U8379 ( .A1(n6422), .A2(n4911), .Y(n8908) );
  NAND2X0_RVT U8380 ( .A1(n8881), .A2(n4961), .Y(n8907) );
  XNOR2X1_RVT U8381 ( .A1(n8909), .A2(n7864), .Y(n8580) );
  NAND2X0_RVT U8382 ( .A1(n8910), .A2(n8911), .Y(n8909) );
  NAND2X0_RVT U8383 ( .A1(n6422), .A2(n4940), .Y(n8911) );
  NAND2X0_RVT U8384 ( .A1(n8881), .A2(n4957), .Y(n8910) );
  XNOR2X1_RVT U8385 ( .A1(n8912), .A2(n7864), .Y(n8594) );
  NAND2X0_RVT U8386 ( .A1(n8913), .A2(n8914), .Y(n8912) );
  NAND2X0_RVT U8387 ( .A1(n6422), .A2(n4941), .Y(n8914) );
  NAND2X0_RVT U8388 ( .A1(n8881), .A2(n4954), .Y(n8913) );
  XNOR2X1_RVT U8389 ( .A1(n8915), .A2(n7864), .Y(n8608) );
  NAND2X0_RVT U8390 ( .A1(n8916), .A2(n8917), .Y(n8915) );
  NAND2X0_RVT U8391 ( .A1(n6422), .A2(n4942), .Y(n8917) );
  NAND2X0_RVT U8392 ( .A1(n8881), .A2(n4956), .Y(n8916) );
  XNOR2X1_RVT U8393 ( .A1(n8918), .A2(n7864), .Y(n8622) );
  NAND2X0_RVT U8394 ( .A1(n8919), .A2(n8920), .Y(n8918) );
  NAND2X0_RVT U8395 ( .A1(n6422), .A2(n4943), .Y(n8920) );
  NAND2X0_RVT U8396 ( .A1(n8881), .A2(n4953), .Y(n8919) );
  XNOR2X1_RVT U8397 ( .A1(n8921), .A2(n7864), .Y(n8636) );
  NAND2X0_RVT U8398 ( .A1(n8922), .A2(n8923), .Y(n8921) );
  NAND2X0_RVT U8399 ( .A1(n6422), .A2(n4966), .Y(n8923) );
  NAND2X0_RVT U8400 ( .A1(n8881), .A2(n4952), .Y(n8922) );
  XNOR2X1_RVT U8401 ( .A1(n8924), .A2(n7864), .Y(n8650) );
  NAND2X0_RVT U8402 ( .A1(n8925), .A2(n8926), .Y(n8924) );
  NAND2X0_RVT U8403 ( .A1(n6422), .A2(n4944), .Y(n8926) );
  NAND2X0_RVT U8404 ( .A1(n8881), .A2(n4955), .Y(n8925) );
  AND2X1_RVT U8405 ( .A1(n9536), .A2(n6422), .Y(n8693) );
  INVX0_RVT U8406 ( .A(n8704), .Y(n8877) );
  NAND2X0_RVT U8407 ( .A1(n9535), .A2(n6422), .Y(n8704) );
  INVX0_RVT U8408 ( .A(n8715), .Y(n8876) );
  NAND2X0_RVT U8409 ( .A1(n9534), .A2(n6422), .Y(n8715) );
  INVX0_RVT U8410 ( .A(n8726), .Y(n8875) );
  NAND2X0_RVT U8411 ( .A1(n9532), .A2(n6422), .Y(n8726) );
  INVX0_RVT U8412 ( .A(n8737), .Y(n8874) );
  NAND2X0_RVT U8413 ( .A1(n9531), .A2(n6422), .Y(n8737) );
  INVX0_RVT U8414 ( .A(n8748), .Y(n8873) );
  NAND2X0_RVT U8415 ( .A1(n9530), .A2(n6422), .Y(n8748) );
  INVX0_RVT U8416 ( .A(n8759), .Y(n8872) );
  NAND2X0_RVT U8417 ( .A1(n9529), .A2(n6422), .Y(n8759) );
  INVX0_RVT U8418 ( .A(n8770), .Y(n8871) );
  NAND2X0_RVT U8419 ( .A1(n9528), .A2(n6422), .Y(n8770) );
  INVX0_RVT U8420 ( .A(n8781), .Y(n8870) );
  NAND2X0_RVT U8421 ( .A1(n9527), .A2(n6422), .Y(n8781) );
  INVX0_RVT U8422 ( .A(n8792), .Y(n8869) );
  NAND2X0_RVT U8423 ( .A1(n9526), .A2(n6422), .Y(n8792) );
  INVX0_RVT U8424 ( .A(n8803), .Y(n8868) );
  NAND2X0_RVT U8425 ( .A1(n9525), .A2(n6422), .Y(n8803) );
  INVX0_RVT U8426 ( .A(n8814), .Y(n8867) );
  NAND2X0_RVT U8427 ( .A1(n9524), .A2(n6422), .Y(n8814) );
  INVX0_RVT U8428 ( .A(n8825), .Y(n8866) );
  NAND2X0_RVT U8429 ( .A1(n9523), .A2(n6422), .Y(n8825) );
  OR2X1_RVT U8430 ( .A1(n6853), .A2(n7910), .Y(n8865) );
  AND2X1_RVT U8431 ( .A1(n9521), .A2(n6422), .Y(n7910) );
  NAND2X0_RVT U8432 ( .A1(n7908), .A2(n7861), .Y(n8929) );
  XNOR2X1_RVT U8433 ( .A1(n8930), .A2(n8931), .Y(n7861) );
  NAND2X0_RVT U8434 ( .A1(n8322), .A2(n8323), .Y(n8931) );
  NAND2X0_RVT U8435 ( .A1(n8932), .A2(n8933), .Y(n8323) );
  NAND2X0_RVT U8436 ( .A1(n8108), .A2(n5056), .Y(n8933) );
  NAND2X0_RVT U8437 ( .A1(rEIP[30]), .A2(n8109), .Y(n8932) );
  AND3X1_RVT U8438 ( .A1(n8317), .A2(n8311), .A3(n8310), .Y(n8322) );
  AND3X1_RVT U8439 ( .A1(n8305), .A2(n8299), .A3(n8298), .Y(n8310) );
  AND3X1_RVT U8440 ( .A1(n8293), .A2(n8287), .A3(n8286), .Y(n8298) );
  AND3X1_RVT U8441 ( .A1(n8281), .A2(n8275), .A3(n8274), .Y(n8286) );
  AND3X1_RVT U8442 ( .A1(n8269), .A2(n8263), .A3(n8262), .Y(n8274) );
  AND3X1_RVT U8443 ( .A1(n8257), .A2(n8251), .A3(n8250), .Y(n8262) );
  AND3X1_RVT U8444 ( .A1(n8245), .A2(n8239), .A3(n8238), .Y(n8250) );
  AND3X1_RVT U8445 ( .A1(n8233), .A2(n8227), .A3(n8226), .Y(n8238) );
  AND3X1_RVT U8446 ( .A1(n8221), .A2(n8215), .A3(n8214), .Y(n8226) );
  AND3X1_RVT U8447 ( .A1(n8209), .A2(n8203), .A3(n8202), .Y(n8214) );
  AND3X1_RVT U8448 ( .A1(n8197), .A2(n8190), .A3(n8189), .Y(n8202) );
  AND2X1_RVT U8449 ( .A1(n8181), .A2(n8180), .Y(n8189) );
  NAND2X0_RVT U8450 ( .A1(n8934), .A2(n8935), .Y(n8180) );
  NAND2X0_RVT U8451 ( .A1(n8108), .A2(n5057), .Y(n8935) );
  NAND2X0_RVT U8452 ( .A1(rEIP[7]), .A2(n8109), .Y(n8934) );
  AND2X1_RVT U8453 ( .A1(n8170), .A2(n8169), .Y(n8181) );
  NAND2X0_RVT U8454 ( .A1(n8936), .A2(n8937), .Y(n8169) );
  NAND2X0_RVT U8455 ( .A1(n8108), .A2(n5058), .Y(n8937) );
  NAND2X0_RVT U8456 ( .A1(rEIP[6]), .A2(n8109), .Y(n8936) );
  AND2X1_RVT U8457 ( .A1(n8159), .A2(n8158), .Y(n8170) );
  NAND2X0_RVT U8458 ( .A1(n8938), .A2(n8939), .Y(n8158) );
  NAND2X0_RVT U8459 ( .A1(n8108), .A2(n5059), .Y(n8939) );
  NAND2X0_RVT U8460 ( .A1(rEIP[5]), .A2(n8109), .Y(n8938) );
  AND2X1_RVT U8461 ( .A1(n8148), .A2(n8147), .Y(n8159) );
  NAND2X0_RVT U8462 ( .A1(n8940), .A2(n8941), .Y(n8147) );
  NAND2X0_RVT U8463 ( .A1(n8108), .A2(n5060), .Y(n8941) );
  NAND2X0_RVT U8464 ( .A1(rEIP[4]), .A2(n8109), .Y(n8940) );
  AND2X1_RVT U8465 ( .A1(n8137), .A2(n8136), .Y(n8148) );
  NAND2X0_RVT U8466 ( .A1(n8942), .A2(n8943), .Y(n8136) );
  NAND2X0_RVT U8467 ( .A1(n8108), .A2(n5061), .Y(n8943) );
  NAND2X0_RVT U8468 ( .A1(rEIP[3]), .A2(n8109), .Y(n8942) );
  AND2X1_RVT U8469 ( .A1(n8944), .A2(n8125), .Y(n8137) );
  NAND2X0_RVT U8470 ( .A1(n8945), .A2(n8946), .Y(n8125) );
  NAND2X0_RVT U8471 ( .A1(n8108), .A2(n5062), .Y(n8946) );
  NAND2X0_RVT U8472 ( .A1(rEIP[2]), .A2(n8109), .Y(n8945) );
  NAND2X0_RVT U8473 ( .A1(n8126), .A2(n8127), .Y(n8944) );
  NAND2X0_RVT U8474 ( .A1(n8118), .A2(n8119), .Y(n8127) );
  NAND2X0_RVT U8475 ( .A1(n8947), .A2(n8948), .Y(n8119) );
  NAND2X0_RVT U8476 ( .A1(n8108), .A2(n5063), .Y(n8948) );
  NAND2X0_RVT U8477 ( .A1(rEIP[1]), .A2(n8109), .Y(n8947) );
  NAND4X0_RVT U8478 ( .A1(n8949), .A2(n8950), .A3(n8951), .A4(n8952), .Y(n8118) );
  NAND2X0_RVT U8479 ( .A1(n8105), .A2(n5128), .Y(n8952) );
  NAND2X0_RVT U8480 ( .A1(n8106), .A2(n8421), .Y(n8951) );
  NAND4X0_RVT U8481 ( .A1(n8953), .A2(n8954), .A3(n8955), .A4(n8956), .Y(n8421) );
  NAND2X0_RVT U8482 ( .A1(n7842), .A2(n8957), .Y(n8956) );
  NAND4X0_RVT U8483 ( .A1(n8958), .A2(n8959), .A3(n8960), .A4(n8961), .Y(n8957) );
  NAND2X0_RVT U8484 ( .A1(n7694), .A2(n5129), .Y(n8961) );
  NAND2X0_RVT U8485 ( .A1(n7678), .A2(n5004), .Y(n8960) );
  NAND2X0_RVT U8486 ( .A1(n7766), .A2(n5005), .Y(n8959) );
  NAND2X0_RVT U8487 ( .A1(n8501), .A2(n5003), .Y(n8958) );
  NAND2X0_RVT U8488 ( .A1(n7853), .A2(n8962), .Y(n8955) );
  NAND2X0_RVT U8489 ( .A1(n7848), .A2(n7742), .Y(n8954) );
  NAND2X0_RVT U8490 ( .A1(n7852), .A2(n7783), .Y(n8953) );
  INVX0_RVT U8491 ( .A(n8109), .Y(n8949) );
  AND3X1_RVT U8492 ( .A1(n8963), .A2(n5390), .A3(n8964), .Y(n8126) );
  NAND2X0_RVT U8493 ( .A1(n8106), .A2(n8417), .Y(n8964) );
  NAND4X0_RVT U8494 ( .A1(n8965), .A2(n8966), .A3(n8967), .A4(n8968), .Y(n8417) );
  NAND2X0_RVT U8495 ( .A1(n7842), .A2(n8969), .Y(n8968) );
  NAND4X0_RVT U8496 ( .A1(n8970), .A2(n8971), .A3(n8972), .A4(n8973), .Y(n8969) );
  NAND2X0_RVT U8497 ( .A1(n7694), .A2(n5130), .Y(n8973) );
  NAND2X0_RVT U8498 ( .A1(n7678), .A2(n5011), .Y(n8972) );
  NAND2X0_RVT U8499 ( .A1(n7766), .A2(n5012), .Y(n8971) );
  NAND2X0_RVT U8500 ( .A1(n8501), .A2(n5010), .Y(n8970) );
  NAND2X0_RVT U8501 ( .A1(n7853), .A2(n8974), .Y(n8967) );
  NAND2X0_RVT U8502 ( .A1(n7848), .A2(n7730), .Y(n8966) );
  NAND2X0_RVT U8503 ( .A1(n7852), .A2(n7793), .Y(n8965) );
  INVX0_RVT U8504 ( .A(n7007), .Y(n8106) );
  NAND2X0_RVT U8505 ( .A1(n8105), .A2(n5131), .Y(n8963) );
  INVX0_RVT U8506 ( .A(n7197), .Y(n8105) );
  NAND3X0_RVT U8507 ( .A1(n8975), .A2(n8976), .A3(n8977), .Y(n8190) );
  NAND2X0_RVT U8508 ( .A1(rEIP[8]), .A2(n8109), .Y(n8977) );
  NAND2X0_RVT U8509 ( .A1(n8978), .A2(n7430), .Y(n8976) );
  NAND4X0_RVT U8510 ( .A1(n8979), .A2(n8980), .A3(n8981), .A4(n8982), .Y(n8978) );
  NAND2X0_RVT U8511 ( .A1(n7848), .A2(n7775), .Y(n8982) );
  NAND3X0_RVT U8512 ( .A1(n8983), .A2(n8984), .A3(n8985), .Y(n7775) );
  NAND2X0_RVT U8513 ( .A1(n7766), .A2(n4996), .Y(n8985) );
  NAND2X0_RVT U8514 ( .A1(n7694), .A2(n4997), .Y(n8984) );
  NAND2X0_RVT U8515 ( .A1(n7678), .A2(n4998), .Y(n8983) );
  NAND2X0_RVT U8516 ( .A1(n7842), .A2(n8502), .Y(n8981) );
  NAND3X0_RVT U8517 ( .A1(n8986), .A2(n8987), .A3(n8988), .Y(n8502) );
  NAND2X0_RVT U8518 ( .A1(n7766), .A2(n4999), .Y(n8988) );
  NAND2X0_RVT U8519 ( .A1(n7694), .A2(n5132), .Y(n8987) );
  NAND2X0_RVT U8520 ( .A1(n7678), .A2(n5000), .Y(n8986) );
  NAND2X0_RVT U8521 ( .A1(n7852), .A2(n7771), .Y(n8980) );
  NAND3X0_RVT U8522 ( .A1(n8989), .A2(n8990), .A3(n8991), .Y(n7771) );
  NAND2X0_RVT U8523 ( .A1(n7766), .A2(n5133), .Y(n8991) );
  NAND2X0_RVT U8524 ( .A1(n7694), .A2(n5134), .Y(n8990) );
  NAND2X0_RVT U8525 ( .A1(n7678), .A2(n5135), .Y(n8989) );
  NAND2X0_RVT U8526 ( .A1(n7853), .A2(n7774), .Y(n8979) );
  NAND3X0_RVT U8527 ( .A1(n8992), .A2(n8993), .A3(n8994), .Y(n7774) );
  NAND2X0_RVT U8528 ( .A1(n7766), .A2(n5001), .Y(n8994) );
  NAND2X0_RVT U8529 ( .A1(n7694), .A2(n5136), .Y(n8993) );
  NAND2X0_RVT U8530 ( .A1(n7678), .A2(n5002), .Y(n8992) );
  NAND2X0_RVT U8531 ( .A1(n8108), .A2(n5064), .Y(n8975) );
  NAND3X0_RVT U8532 ( .A1(n8995), .A2(n8996), .A3(n8997), .Y(n8197) );
  NAND2X0_RVT U8533 ( .A1(rEIP[9]), .A2(n8109), .Y(n8997) );
  NAND2X0_RVT U8534 ( .A1(n8998), .A2(n7430), .Y(n8996) );
  NAND4X0_RVT U8535 ( .A1(n8999), .A2(n9000), .A3(n9001), .A4(n9002), .Y(n8998) );
  NAND2X0_RVT U8536 ( .A1(n7848), .A2(n7744), .Y(n9002) );
  NAND3X0_RVT U8537 ( .A1(n9003), .A2(n9004), .A3(n9005), .Y(n7744) );
  NAND2X0_RVT U8538 ( .A1(n7766), .A2(n5003), .Y(n9005) );
  NAND2X0_RVT U8539 ( .A1(n7694), .A2(n5004), .Y(n9004) );
  NAND2X0_RVT U8540 ( .A1(n7678), .A2(n5005), .Y(n9003) );
  NAND2X0_RVT U8541 ( .A1(n7842), .A2(n8962), .Y(n9001) );
  NAND3X0_RVT U8542 ( .A1(n9006), .A2(n9007), .A3(n9008), .Y(n8962) );
  NAND2X0_RVT U8543 ( .A1(n7766), .A2(n5006), .Y(n9008) );
  NAND2X0_RVT U8544 ( .A1(n7694), .A2(n5137), .Y(n9007) );
  NAND2X0_RVT U8545 ( .A1(n7678), .A2(n5007), .Y(n9006) );
  NAND2X0_RVT U8546 ( .A1(n7852), .A2(n7742), .Y(n9000) );
  NAND3X0_RVT U8547 ( .A1(n9009), .A2(n9010), .A3(n9011), .Y(n7742) );
  NAND2X0_RVT U8548 ( .A1(n7766), .A2(n5138), .Y(n9011) );
  NAND2X0_RVT U8549 ( .A1(n7694), .A2(n5139), .Y(n9010) );
  NAND2X0_RVT U8550 ( .A1(n7678), .A2(n5140), .Y(n9009) );
  NAND2X0_RVT U8551 ( .A1(n7853), .A2(n7783), .Y(n8999) );
  NAND3X0_RVT U8552 ( .A1(n9012), .A2(n9013), .A3(n9014), .Y(n7783) );
  NAND2X0_RVT U8553 ( .A1(n7766), .A2(n5008), .Y(n9014) );
  NAND2X0_RVT U8554 ( .A1(n7694), .A2(n5141), .Y(n9013) );
  NAND2X0_RVT U8555 ( .A1(n7678), .A2(n5009), .Y(n9012) );
  NAND2X0_RVT U8556 ( .A1(n8108), .A2(n5065), .Y(n8995) );
  NAND3X0_RVT U8557 ( .A1(n9015), .A2(n9016), .A3(n9017), .Y(n8203) );
  NAND2X0_RVT U8558 ( .A1(rEIP[10]), .A2(n8109), .Y(n9017) );
  NAND2X0_RVT U8559 ( .A1(n9018), .A2(n7430), .Y(n9016) );
  NAND4X0_RVT U8560 ( .A1(n9019), .A2(n9020), .A3(n9021), .A4(n9022), .Y(n9018) );
  NAND2X0_RVT U8561 ( .A1(n7848), .A2(n7732), .Y(n9022) );
  NAND3X0_RVT U8562 ( .A1(n9023), .A2(n9024), .A3(n9025), .Y(n7732) );
  NAND2X0_RVT U8563 ( .A1(n7766), .A2(n5010), .Y(n9025) );
  NAND2X0_RVT U8564 ( .A1(n7694), .A2(n5011), .Y(n9024) );
  NAND2X0_RVT U8565 ( .A1(n7678), .A2(n5012), .Y(n9023) );
  NAND2X0_RVT U8566 ( .A1(n7842), .A2(n8974), .Y(n9021) );
  NAND3X0_RVT U8567 ( .A1(n9026), .A2(n9027), .A3(n9028), .Y(n8974) );
  NAND2X0_RVT U8568 ( .A1(n7766), .A2(n5013), .Y(n9028) );
  NAND2X0_RVT U8569 ( .A1(n7694), .A2(n5142), .Y(n9027) );
  NAND2X0_RVT U8570 ( .A1(n7678), .A2(n5014), .Y(n9026) );
  NAND2X0_RVT U8571 ( .A1(n7852), .A2(n7730), .Y(n9020) );
  NAND3X0_RVT U8572 ( .A1(n9029), .A2(n9030), .A3(n9031), .Y(n7730) );
  NAND2X0_RVT U8573 ( .A1(n7766), .A2(n5143), .Y(n9031) );
  NAND2X0_RVT U8574 ( .A1(n7694), .A2(n5144), .Y(n9030) );
  NAND2X0_RVT U8575 ( .A1(n7678), .A2(n5145), .Y(n9029) );
  NAND2X0_RVT U8576 ( .A1(n7853), .A2(n7793), .Y(n9019) );
  NAND3X0_RVT U8577 ( .A1(n9032), .A2(n9033), .A3(n9034), .Y(n7793) );
  NAND2X0_RVT U8578 ( .A1(n7766), .A2(n5015), .Y(n9034) );
  NAND2X0_RVT U8579 ( .A1(n7694), .A2(n5146), .Y(n9033) );
  NAND2X0_RVT U8580 ( .A1(n7678), .A2(n5108), .Y(n9032) );
  NAND2X0_RVT U8581 ( .A1(n8108), .A2(n5066), .Y(n9015) );
  NAND3X0_RVT U8582 ( .A1(n9035), .A2(n9036), .A3(n9037), .Y(n8209) );
  NAND2X0_RVT U8583 ( .A1(rEIP[11]), .A2(n8109), .Y(n9037) );
  NAND2X0_RVT U8584 ( .A1(n9038), .A2(n7430), .Y(n9036) );
  NAND4X0_RVT U8585 ( .A1(n9039), .A2(n9040), .A3(n9041), .A4(n9042), .Y(n9038) );
  NAND2X0_RVT U8586 ( .A1(n7848), .A2(n7721), .Y(n9042) );
  NAND3X0_RVT U8587 ( .A1(n9043), .A2(n9044), .A3(n9045), .Y(n7721) );
  NAND2X0_RVT U8588 ( .A1(n7766), .A2(n5016), .Y(n9045) );
  NAND2X0_RVT U8589 ( .A1(n7694), .A2(n5017), .Y(n9044) );
  NAND2X0_RVT U8590 ( .A1(n7678), .A2(n5018), .Y(n9043) );
  NAND2X0_RVT U8591 ( .A1(n7842), .A2(n8527), .Y(n9041) );
  NAND3X0_RVT U8592 ( .A1(n9046), .A2(n9047), .A3(n9048), .Y(n8527) );
  NAND2X0_RVT U8593 ( .A1(n7766), .A2(n5019), .Y(n9048) );
  NAND2X0_RVT U8594 ( .A1(n7694), .A2(n5147), .Y(n9047) );
  NAND2X0_RVT U8595 ( .A1(n7678), .A2(n5020), .Y(n9046) );
  NAND2X0_RVT U8596 ( .A1(n7852), .A2(n7719), .Y(n9040) );
  NAND3X0_RVT U8597 ( .A1(n9049), .A2(n9050), .A3(n9051), .Y(n7719) );
  NAND2X0_RVT U8598 ( .A1(n7766), .A2(n5148), .Y(n9051) );
  NAND2X0_RVT U8599 ( .A1(n7694), .A2(n5149), .Y(n9050) );
  NAND2X0_RVT U8600 ( .A1(n7678), .A2(n5150), .Y(n9049) );
  NAND2X0_RVT U8601 ( .A1(n7853), .A2(n7803), .Y(n9039) );
  NAND3X0_RVT U8602 ( .A1(n9052), .A2(n9053), .A3(n9054), .Y(n7803) );
  NAND2X0_RVT U8603 ( .A1(n7766), .A2(n5021), .Y(n9054) );
  NAND2X0_RVT U8604 ( .A1(n7694), .A2(n5151), .Y(n9053) );
  NAND2X0_RVT U8605 ( .A1(n7678), .A2(n5022), .Y(n9052) );
  NAND2X0_RVT U8606 ( .A1(n8108), .A2(n5067), .Y(n9035) );
  NAND3X0_RVT U8607 ( .A1(n9055), .A2(n9056), .A3(n9057), .Y(n8215) );
  NAND2X0_RVT U8608 ( .A1(rEIP[12]), .A2(n8109), .Y(n9057) );
  NAND2X0_RVT U8609 ( .A1(n9058), .A2(n7430), .Y(n9056) );
  NAND4X0_RVT U8610 ( .A1(n9059), .A2(n9060), .A3(n9061), .A4(n9062), .Y(n9058) );
  NAND2X0_RVT U8611 ( .A1(n7848), .A2(n7709), .Y(n9062) );
  NAND3X0_RVT U8612 ( .A1(n9063), .A2(n9064), .A3(n9065), .Y(n7709) );
  NAND2X0_RVT U8613 ( .A1(n7766), .A2(n5023), .Y(n9065) );
  NAND2X0_RVT U8614 ( .A1(n7694), .A2(n5024), .Y(n9064) );
  NAND2X0_RVT U8615 ( .A1(n7678), .A2(n5025), .Y(n9063) );
  NAND2X0_RVT U8616 ( .A1(n7842), .A2(n8537), .Y(n9061) );
  NAND3X0_RVT U8617 ( .A1(n9066), .A2(n9067), .A3(n9068), .Y(n8537) );
  NAND2X0_RVT U8618 ( .A1(n7766), .A2(n5026), .Y(n9068) );
  NAND2X0_RVT U8619 ( .A1(n7694), .A2(n5152), .Y(n9067) );
  NAND2X0_RVT U8620 ( .A1(n7678), .A2(n5027), .Y(n9066) );
  NAND2X0_RVT U8621 ( .A1(n7852), .A2(n7707), .Y(n9060) );
  NAND3X0_RVT U8622 ( .A1(n9069), .A2(n9070), .A3(n9071), .Y(n7707) );
  NAND2X0_RVT U8623 ( .A1(n7766), .A2(n5153), .Y(n9071) );
  NAND2X0_RVT U8624 ( .A1(n7694), .A2(n5154), .Y(n9070) );
  NAND2X0_RVT U8625 ( .A1(n7678), .A2(n5155), .Y(n9069) );
  NAND2X0_RVT U8626 ( .A1(n7853), .A2(n7813), .Y(n9059) );
  NAND3X0_RVT U8627 ( .A1(n9072), .A2(n9073), .A3(n9074), .Y(n7813) );
  NAND2X0_RVT U8628 ( .A1(n7766), .A2(n5028), .Y(n9074) );
  NAND2X0_RVT U8629 ( .A1(n7694), .A2(n5156), .Y(n9073) );
  NAND2X0_RVT U8630 ( .A1(n7678), .A2(n5029), .Y(n9072) );
  NAND2X0_RVT U8631 ( .A1(n8108), .A2(n5068), .Y(n9055) );
  NAND3X0_RVT U8632 ( .A1(n9075), .A2(n9076), .A3(n9077), .Y(n8221) );
  NAND2X0_RVT U8633 ( .A1(rEIP[13]), .A2(n8109), .Y(n9077) );
  NAND2X0_RVT U8634 ( .A1(n9078), .A2(n7430), .Y(n9076) );
  NAND4X0_RVT U8635 ( .A1(n9079), .A2(n9080), .A3(n9081), .A4(n9082), .Y(n9078) );
  NAND2X0_RVT U8636 ( .A1(n7848), .A2(n7697), .Y(n9082) );
  NAND3X0_RVT U8637 ( .A1(n9083), .A2(n9084), .A3(n9085), .Y(n7697) );
  NAND2X0_RVT U8638 ( .A1(n7766), .A2(n5030), .Y(n9085) );
  NAND2X0_RVT U8639 ( .A1(n7694), .A2(n5031), .Y(n9084) );
  NAND2X0_RVT U8640 ( .A1(n7678), .A2(n5032), .Y(n9083) );
  NAND2X0_RVT U8641 ( .A1(n7842), .A2(n8547), .Y(n9081) );
  NAND3X0_RVT U8642 ( .A1(n9086), .A2(n9087), .A3(n9088), .Y(n8547) );
  NAND2X0_RVT U8643 ( .A1(n7766), .A2(n5033), .Y(n9088) );
  NAND2X0_RVT U8644 ( .A1(n7694), .A2(n5157), .Y(n9087) );
  NAND2X0_RVT U8645 ( .A1(n7678), .A2(n5034), .Y(n9086) );
  NAND2X0_RVT U8646 ( .A1(n7852), .A2(n7695), .Y(n9080) );
  NAND3X0_RVT U8647 ( .A1(n9089), .A2(n9090), .A3(n9091), .Y(n7695) );
  NAND2X0_RVT U8648 ( .A1(n7766), .A2(n5158), .Y(n9091) );
  NAND2X0_RVT U8649 ( .A1(n7694), .A2(n5159), .Y(n9090) );
  NAND2X0_RVT U8650 ( .A1(n7678), .A2(n5160), .Y(n9089) );
  NAND2X0_RVT U8651 ( .A1(n7853), .A2(n7823), .Y(n9079) );
  NAND3X0_RVT U8652 ( .A1(n9092), .A2(n9093), .A3(n9094), .Y(n7823) );
  NAND2X0_RVT U8653 ( .A1(n7766), .A2(n5035), .Y(n9094) );
  NAND2X0_RVT U8654 ( .A1(n7694), .A2(n5161), .Y(n9093) );
  NAND2X0_RVT U8655 ( .A1(n7678), .A2(n5036), .Y(n9092) );
  NAND2X0_RVT U8656 ( .A1(n8108), .A2(n5069), .Y(n9075) );
  NAND3X0_RVT U8657 ( .A1(n9095), .A2(n9096), .A3(n9097), .Y(n8227) );
  NAND2X0_RVT U8658 ( .A1(rEIP[14]), .A2(n8109), .Y(n9097) );
  NAND2X0_RVT U8659 ( .A1(n9098), .A2(n7430), .Y(n9096) );
  NAND4X0_RVT U8660 ( .A1(n9099), .A2(n9100), .A3(n9101), .A4(n9102), .Y(n9098) );
  NAND2X0_RVT U8661 ( .A1(n7848), .A2(n7684), .Y(n9102) );
  NAND3X0_RVT U8662 ( .A1(n9103), .A2(n9104), .A3(n9105), .Y(n7684) );
  NAND2X0_RVT U8663 ( .A1(n7766), .A2(n5037), .Y(n9105) );
  NAND2X0_RVT U8664 ( .A1(n7694), .A2(n5038), .Y(n9104) );
  NAND2X0_RVT U8665 ( .A1(n7678), .A2(n5039), .Y(n9103) );
  NAND2X0_RVT U8666 ( .A1(n7842), .A2(n8557), .Y(n9101) );
  NAND3X0_RVT U8667 ( .A1(n9106), .A2(n9107), .A3(n9108), .Y(n8557) );
  NAND2X0_RVT U8668 ( .A1(n7766), .A2(n5040), .Y(n9108) );
  NAND2X0_RVT U8669 ( .A1(n7694), .A2(n5162), .Y(n9107) );
  NAND2X0_RVT U8670 ( .A1(n7678), .A2(n5041), .Y(n9106) );
  NAND2X0_RVT U8671 ( .A1(n7852), .A2(n7680), .Y(n9100) );
  NAND3X0_RVT U8672 ( .A1(n9109), .A2(n9110), .A3(n9111), .Y(n7680) );
  NAND2X0_RVT U8673 ( .A1(n7766), .A2(n5163), .Y(n9111) );
  NAND2X0_RVT U8674 ( .A1(n7694), .A2(n5164), .Y(n9110) );
  NAND2X0_RVT U8675 ( .A1(n7678), .A2(n5165), .Y(n9109) );
  NAND2X0_RVT U8676 ( .A1(n7853), .A2(n7762), .Y(n9099) );
  NAND3X0_RVT U8677 ( .A1(n9112), .A2(n9113), .A3(n9114), .Y(n7762) );
  NAND2X0_RVT U8678 ( .A1(n7766), .A2(n5042), .Y(n9114) );
  NAND2X0_RVT U8679 ( .A1(n7694), .A2(n5166), .Y(n9113) );
  NAND2X0_RVT U8680 ( .A1(n7678), .A2(n5109), .Y(n9112) );
  NAND2X0_RVT U8681 ( .A1(n8108), .A2(n5070), .Y(n9095) );
  NAND3X0_RVT U8682 ( .A1(n9115), .A2(n9116), .A3(n9117), .Y(n8233) );
  NAND2X0_RVT U8683 ( .A1(rEIP[15]), .A2(n8109), .Y(n9117) );
  NAND2X0_RVT U8684 ( .A1(n9118), .A2(n7430), .Y(n9116) );
  NAND2X0_RVT U8685 ( .A1(n9119), .A2(n7009), .Y(n7197) );
  INVX0_RVT U8686 ( .A(n6727), .Y(n9119) );
  NAND2X0_RVT U8687 ( .A1(n9120), .A2(n7009), .Y(n7007) );
  INVX0_RVT U8688 ( .A(n9121), .Y(n9120) );
  NAND4X0_RVT U8689 ( .A1(n9122), .A2(n9123), .A3(n9124), .A4(n9125), .Y(n9118) );
  NAND2X0_RVT U8690 ( .A1(n7848), .A2(n7754), .Y(n9125) );
  NAND3X0_RVT U8691 ( .A1(n9126), .A2(n9127), .A3(n9128), .Y(n7754) );
  NAND2X0_RVT U8692 ( .A1(n7766), .A2(n5045), .Y(n9128) );
  NAND2X0_RVT U8693 ( .A1(n7694), .A2(n5043), .Y(n9127) );
  NAND2X0_RVT U8694 ( .A1(n7678), .A2(n5044), .Y(n9126) );
  NAND2X0_RVT U8695 ( .A1(n7842), .A2(n9129), .Y(n9124) );
  NAND2X0_RVT U8696 ( .A1(n7852), .A2(n7750), .Y(n9123) );
  NAND2X0_RVT U8697 ( .A1(n7853), .A2(n7753), .Y(n9122) );
  NAND2X0_RVT U8698 ( .A1(n8108), .A2(n5071), .Y(n9115) );
  NAND2X0_RVT U8699 ( .A1(n9130), .A2(n9131), .Y(n8239) );
  NAND2X0_RVT U8700 ( .A1(n8108), .A2(n5072), .Y(n9131) );
  NAND2X0_RVT U8701 ( .A1(rEIP[16]), .A2(n8109), .Y(n9130) );
  NAND2X0_RVT U8702 ( .A1(n9132), .A2(n9133), .Y(n8245) );
  NAND2X0_RVT U8703 ( .A1(n8108), .A2(n5073), .Y(n9133) );
  NAND2X0_RVT U8704 ( .A1(rEIP[17]), .A2(n8109), .Y(n9132) );
  NAND2X0_RVT U8705 ( .A1(n9134), .A2(n9135), .Y(n8251) );
  NAND2X0_RVT U8706 ( .A1(n8108), .A2(n5074), .Y(n9135) );
  NAND2X0_RVT U8707 ( .A1(rEIP[18]), .A2(n8109), .Y(n9134) );
  NAND2X0_RVT U8708 ( .A1(n9136), .A2(n9137), .Y(n8257) );
  NAND2X0_RVT U8709 ( .A1(n8108), .A2(n5075), .Y(n9137) );
  NAND2X0_RVT U8710 ( .A1(rEIP[19]), .A2(n8109), .Y(n9136) );
  NAND2X0_RVT U8711 ( .A1(n9138), .A2(n9139), .Y(n8263) );
  NAND2X0_RVT U8712 ( .A1(n8108), .A2(n5076), .Y(n9139) );
  NAND2X0_RVT U8713 ( .A1(rEIP[20]), .A2(n8109), .Y(n9138) );
  NAND2X0_RVT U8714 ( .A1(n9140), .A2(n9141), .Y(n8269) );
  NAND2X0_RVT U8715 ( .A1(n8108), .A2(n5077), .Y(n9141) );
  NAND2X0_RVT U8716 ( .A1(rEIP[21]), .A2(n8109), .Y(n9140) );
  NAND2X0_RVT U8717 ( .A1(n9142), .A2(n9143), .Y(n8275) );
  NAND2X0_RVT U8718 ( .A1(n8108), .A2(n5078), .Y(n9143) );
  NAND2X0_RVT U8719 ( .A1(rEIP[22]), .A2(n8109), .Y(n9142) );
  NAND2X0_RVT U8720 ( .A1(n9144), .A2(n9145), .Y(n8281) );
  NAND2X0_RVT U8721 ( .A1(n8108), .A2(n5079), .Y(n9145) );
  NAND2X0_RVT U8722 ( .A1(rEIP[23]), .A2(n8109), .Y(n9144) );
  NAND2X0_RVT U8723 ( .A1(n9146), .A2(n9147), .Y(n8287) );
  NAND2X0_RVT U8724 ( .A1(n8108), .A2(n5080), .Y(n9147) );
  NAND2X0_RVT U8725 ( .A1(rEIP[24]), .A2(n8109), .Y(n9146) );
  NAND2X0_RVT U8726 ( .A1(n9148), .A2(n9149), .Y(n8293) );
  NAND2X0_RVT U8727 ( .A1(n8108), .A2(n5081), .Y(n9149) );
  NAND2X0_RVT U8728 ( .A1(rEIP[25]), .A2(n8109), .Y(n9148) );
  NAND2X0_RVT U8729 ( .A1(n9150), .A2(n9151), .Y(n8299) );
  NAND2X0_RVT U8730 ( .A1(n8108), .A2(n5082), .Y(n9151) );
  NAND2X0_RVT U8731 ( .A1(rEIP[26]), .A2(n8109), .Y(n9150) );
  NAND2X0_RVT U8732 ( .A1(n9152), .A2(n9153), .Y(n8305) );
  NAND2X0_RVT U8733 ( .A1(n8108), .A2(n5083), .Y(n9153) );
  NAND2X0_RVT U8734 ( .A1(rEIP[27]), .A2(n8109), .Y(n9152) );
  NAND2X0_RVT U8735 ( .A1(n9154), .A2(n9155), .Y(n8311) );
  NAND2X0_RVT U8736 ( .A1(n8108), .A2(n5084), .Y(n9155) );
  NAND2X0_RVT U8737 ( .A1(rEIP[28]), .A2(n8109), .Y(n9154) );
  NAND2X0_RVT U8738 ( .A1(n9156), .A2(n9157), .Y(n8317) );
  NAND2X0_RVT U8739 ( .A1(n8108), .A2(n5085), .Y(n9157) );
  NAND2X0_RVT U8740 ( .A1(rEIP[29]), .A2(n8109), .Y(n9156) );
  NAND2X0_RVT U8741 ( .A1(n9158), .A2(n9159), .Y(n8930) );
  NAND2X0_RVT U8742 ( .A1(n8108), .A2(n5086), .Y(n9159) );
  NAND2X0_RVT U8743 ( .A1(n5371), .A2(n4967), .Y(n5390) );
  INVX0_RVT U8744 ( .A(n6308), .Y(n8950) );
  NAND2X0_RVT U8745 ( .A1(n6531), .A2(n5368), .Y(n6308) );
  NAND3X0_RVT U8746 ( .A1(n791), .A2(n4905), .A3(n8560), .Y(n5368) );
  NAND2X0_RVT U8747 ( .A1(rEIP[31]), .A2(n8109), .Y(n9158) );
  NAND2X0_RVT U8748 ( .A1(n7875), .A2(n755), .Y(n9160) );
  INVX0_RVT U8749 ( .A(n7008), .Y(n7875) );
  NAND3X0_RVT U8750 ( .A1(n7009), .A2(n5268), .A3(n7046), .Y(n7008) );
  INVX0_RVT U8751 ( .A(n7869), .Y(n7871) );
  NAND2X0_RVT U8752 ( .A1(n755), .A2(n5268), .Y(n7869) );
  INVX0_RVT U8753 ( .A(READY_n), .Y(n5268) );
  INVX0_RVT U8754 ( .A(n6531), .Y(n7908) );
  NAND2X0_RVT U8755 ( .A1(n755), .A2(n5371), .Y(n6531) );
  NAND3X0_RVT U8756 ( .A1(n790), .A2(n4910), .A3(n8560), .Y(n5351) );
  NAND3X0_RVT U8757 ( .A1(n7009), .A2(n4958), .A3(n7046), .Y(n8928) );
  INVX0_RVT U8758 ( .A(n8511), .Y(n7046) );
  OR2X1_RVT U8759 ( .A1(n5382), .A2(n9567), .Y(n8927) );
  NAND2X0_RVT U8760 ( .A1(n5357), .A2(n5110), .Y(n5382) );
  INVX0_RVT U8761 ( .A(n5339), .Y(n5357) );
  NAND3X0_RVT U8762 ( .A1(n4905), .A2(n4910), .A3(n6534), .Y(n5339) );
  XOR2X1_RVT U8763 ( .A1(n9161), .A2(n8863), .Y(n6853) );
  NAND2X0_RVT U8764 ( .A1(n9162), .A2(n9163), .Y(n8863) );
  NAND2X0_RVT U8765 ( .A1(n8826), .A2(n8828), .Y(n9163) );
  AND2X1_RVT U8766 ( .A1(n5207), .A2(n4949), .Y(n8826) );
  NAND2X0_RVT U8767 ( .A1(n8827), .A2(n8828), .Y(n9162) );
  NAND2X0_RVT U8768 ( .A1(n9164), .A2(n9165), .Y(n8828) );
  NAND2X0_RVT U8769 ( .A1(n8815), .A2(n8817), .Y(n9165) );
  AND2X1_RVT U8770 ( .A1(n5206), .A2(n4955), .Y(n8815) );
  NAND2X0_RVT U8771 ( .A1(n8816), .A2(n8817), .Y(n9164) );
  NAND2X0_RVT U8772 ( .A1(n9166), .A2(n9167), .Y(n8817) );
  NAND2X0_RVT U8773 ( .A1(n8804), .A2(n8806), .Y(n9167) );
  AND2X1_RVT U8774 ( .A1(n5205), .A2(n4946), .Y(n8804) );
  NAND2X0_RVT U8775 ( .A1(n8805), .A2(n8806), .Y(n9166) );
  NAND2X0_RVT U8776 ( .A1(n9168), .A2(n9169), .Y(n8806) );
  NAND2X0_RVT U8777 ( .A1(n8793), .A2(n8795), .Y(n9169) );
  AND2X1_RVT U8778 ( .A1(n5204), .A2(n4952), .Y(n8793) );
  NAND2X0_RVT U8779 ( .A1(n8794), .A2(n8795), .Y(n9168) );
  NAND2X0_RVT U8780 ( .A1(n9170), .A2(n9171), .Y(n8795) );
  NAND2X0_RVT U8781 ( .A1(n8782), .A2(n8784), .Y(n9171) );
  AND2X1_RVT U8782 ( .A1(n5207), .A2(n4947), .Y(n8782) );
  NAND2X0_RVT U8783 ( .A1(n8783), .A2(n8784), .Y(n9170) );
  NAND2X0_RVT U8784 ( .A1(n9172), .A2(n9173), .Y(n8784) );
  NAND2X0_RVT U8785 ( .A1(n8771), .A2(n8773), .Y(n9173) );
  AND2X1_RVT U8786 ( .A1(n5206), .A2(n4953), .Y(n8771) );
  NAND2X0_RVT U8787 ( .A1(n8772), .A2(n8773), .Y(n9172) );
  NAND2X0_RVT U8788 ( .A1(n9174), .A2(n9175), .Y(n8773) );
  NAND2X0_RVT U8789 ( .A1(n8760), .A2(n8762), .Y(n9175) );
  AND2X1_RVT U8790 ( .A1(n5205), .A2(n4950), .Y(n8760) );
  NAND2X0_RVT U8791 ( .A1(n8761), .A2(n8762), .Y(n9174) );
  NAND2X0_RVT U8792 ( .A1(n9176), .A2(n9177), .Y(n8762) );
  NAND2X0_RVT U8793 ( .A1(n8749), .A2(n8751), .Y(n9177) );
  AND2X1_RVT U8794 ( .A1(n5204), .A2(n4956), .Y(n8749) );
  NAND2X0_RVT U8795 ( .A1(n8750), .A2(n8751), .Y(n9176) );
  NAND2X0_RVT U8796 ( .A1(n9178), .A2(n9179), .Y(n8751) );
  NAND2X0_RVT U8797 ( .A1(n8738), .A2(n8740), .Y(n9179) );
  AND2X1_RVT U8798 ( .A1(n5207), .A2(n4948), .Y(n8738) );
  NAND2X0_RVT U8799 ( .A1(n8739), .A2(n8740), .Y(n9178) );
  NAND2X0_RVT U8800 ( .A1(n9180), .A2(n9181), .Y(n8740) );
  NAND2X0_RVT U8801 ( .A1(n8727), .A2(n8729), .Y(n9181) );
  AND2X1_RVT U8802 ( .A1(n5206), .A2(n4954), .Y(n8727) );
  NAND2X0_RVT U8803 ( .A1(n8728), .A2(n8729), .Y(n9180) );
  NAND2X0_RVT U8804 ( .A1(n9182), .A2(n9183), .Y(n8729) );
  NAND2X0_RVT U8805 ( .A1(n8716), .A2(n8718), .Y(n9183) );
  AND2X1_RVT U8806 ( .A1(n5205), .A2(n4951), .Y(n8716) );
  NAND2X0_RVT U8807 ( .A1(n8717), .A2(n8718), .Y(n9182) );
  NAND2X0_RVT U8808 ( .A1(n9184), .A2(n9185), .Y(n8718) );
  NAND2X0_RVT U8809 ( .A1(n8705), .A2(n8707), .Y(n9185) );
  AND2X1_RVT U8810 ( .A1(n5204), .A2(n4957), .Y(n8705) );
  NAND2X0_RVT U8811 ( .A1(n8706), .A2(n8707), .Y(n9184) );
  NAND2X0_RVT U8812 ( .A1(n9186), .A2(n9187), .Y(n8707) );
  OR2X1_RVT U8813 ( .A1(n9188), .A2(n8694), .Y(n9187) );
  NAND2X0_RVT U8814 ( .A1(n5207), .A2(n4959), .Y(n8694) );
  NAND2X0_RVT U8815 ( .A1(n8696), .A2(n8695), .Y(n9186) );
  NAND2X0_RVT U8816 ( .A1(n9189), .A2(n9190), .Y(n8695) );
  NAND2X0_RVT U8817 ( .A1(n5214), .A2(n5175), .Y(n9190) );
  NAND2X0_RVT U8818 ( .A1(n9191), .A2(n5087), .Y(n9189) );
  INVX0_RVT U8819 ( .A(n9188), .Y(n8696) );
  NAND2X0_RVT U8820 ( .A1(n8685), .A2(n8684), .Y(n9188) );
  NAND2X0_RVT U8821 ( .A1(n9192), .A2(n9193), .Y(n8684) );
  NAND2X0_RVT U8822 ( .A1(n5206), .A2(n4961), .Y(n9193) );
  NAND3X0_RVT U8823 ( .A1(n9194), .A2(n5054), .A3(n9191), .Y(n9192) );
  OR4X1_RVT U8824 ( .A1(n9195), .A2(n9196), .A3(n9197), .A4(n9198), .Y(n9194)
         );
  NAND4X0_RVT U8825 ( .A1(n9553), .A2(n9554), .A3(n9555), .A4(n9556), .Y(n9198) );
  NAND4X0_RVT U8826 ( .A1(n9557), .A2(n9558), .A3(n9559), .A4(n9560), .Y(n9197) );
  NAND4X0_RVT U8827 ( .A1(n9545), .A2(n9546), .A3(n9547), .A4(n9548), .Y(n9196) );
  NAND4X0_RVT U8828 ( .A1(n9549), .A2(n9550), .A3(n9551), .A4(n9552), .Y(n9195) );
  NAND3X0_RVT U8829 ( .A1(n9199), .A2(n7006), .A3(n9200), .Y(n8685) );
  NAND2X0_RVT U8830 ( .A1(n9191), .A2(n5088), .Y(n9200) );
  NAND2X0_RVT U8831 ( .A1(n5213), .A2(n5176), .Y(n9199) );
  NAND2X0_RVT U8832 ( .A1(n9201), .A2(n9202), .Y(n8706) );
  NAND2X0_RVT U8833 ( .A1(n5212), .A2(n5177), .Y(n9202) );
  NAND2X0_RVT U8834 ( .A1(n9191), .A2(n5089), .Y(n9201) );
  NAND2X0_RVT U8835 ( .A1(n9203), .A2(n9204), .Y(n8717) );
  NAND2X0_RVT U8836 ( .A1(n5215), .A2(n5178), .Y(n9204) );
  NAND2X0_RVT U8837 ( .A1(n9191), .A2(n5090), .Y(n9203) );
  NAND2X0_RVT U8838 ( .A1(n9205), .A2(n9206), .Y(n8728) );
  NAND2X0_RVT U8839 ( .A1(n5214), .A2(n5179), .Y(n9206) );
  NAND2X0_RVT U8840 ( .A1(n9191), .A2(n5091), .Y(n9205) );
  NAND2X0_RVT U8841 ( .A1(n9207), .A2(n9208), .Y(n8739) );
  NAND2X0_RVT U8842 ( .A1(n5213), .A2(n5180), .Y(n9208) );
  NAND2X0_RVT U8843 ( .A1(n9191), .A2(n5092), .Y(n9207) );
  NAND2X0_RVT U8844 ( .A1(n9209), .A2(n9210), .Y(n8750) );
  NAND2X0_RVT U8845 ( .A1(n5212), .A2(n5181), .Y(n9210) );
  NAND2X0_RVT U8846 ( .A1(n9191), .A2(n5093), .Y(n9209) );
  NAND2X0_RVT U8847 ( .A1(n9211), .A2(n9212), .Y(n8761) );
  NAND2X0_RVT U8848 ( .A1(n5215), .A2(n5182), .Y(n9212) );
  NAND2X0_RVT U8849 ( .A1(n9191), .A2(n5094), .Y(n9211) );
  NAND2X0_RVT U8850 ( .A1(n9213), .A2(n9214), .Y(n8772) );
  NAND2X0_RVT U8851 ( .A1(n5214), .A2(n5183), .Y(n9214) );
  NAND2X0_RVT U8852 ( .A1(n9191), .A2(n5095), .Y(n9213) );
  NAND2X0_RVT U8853 ( .A1(n9215), .A2(n9216), .Y(n8783) );
  NAND2X0_RVT U8854 ( .A1(n5213), .A2(n5184), .Y(n9216) );
  NAND2X0_RVT U8855 ( .A1(n9191), .A2(n5096), .Y(n9215) );
  NAND2X0_RVT U8856 ( .A1(n9217), .A2(n9218), .Y(n8794) );
  NAND2X0_RVT U8857 ( .A1(n5212), .A2(n5185), .Y(n9218) );
  NAND2X0_RVT U8858 ( .A1(n9191), .A2(n5097), .Y(n9217) );
  NAND2X0_RVT U8859 ( .A1(n9219), .A2(n9220), .Y(n8805) );
  NAND2X0_RVT U8860 ( .A1(n5215), .A2(n5186), .Y(n9220) );
  NAND2X0_RVT U8861 ( .A1(n9191), .A2(n5098), .Y(n9219) );
  NAND2X0_RVT U8862 ( .A1(n9221), .A2(n9222), .Y(n8816) );
  NAND2X0_RVT U8863 ( .A1(n5214), .A2(n5187), .Y(n9222) );
  NAND2X0_RVT U8864 ( .A1(n9191), .A2(n5099), .Y(n9221) );
  NAND2X0_RVT U8865 ( .A1(n9223), .A2(n9224), .Y(n8827) );
  NAND2X0_RVT U8866 ( .A1(n5213), .A2(n5188), .Y(n9224) );
  NAND2X0_RVT U8867 ( .A1(n9191), .A2(n5100), .Y(n9223) );
  NAND3X0_RVT U8868 ( .A1(n9225), .A2(n8864), .A3(n9226), .Y(n9161) );
  NAND2X0_RVT U8869 ( .A1(n5212), .A2(n5189), .Y(n9226) );
  NAND2X0_RVT U8870 ( .A1(n5205), .A2(n4960), .Y(n8864) );
  NAND4X0_RVT U8871 ( .A1(n8512), .A2(n7844), .A3(n8514), .A4(n5265), .Y(n7006) );
  AND3X1_RVT U8872 ( .A1(n9227), .A2(n8513), .A3(n9228), .Y(n7844) );
  AND4X1_RVT U8873 ( .A1(n9229), .A2(n9230), .A3(n9231), .A4(n6387), .Y(n8513)
         );
  NAND2X0_RVT U8874 ( .A1(n9191), .A2(n5101), .Y(n9225) );
  INVX0_RVT U8875 ( .A(n7047), .Y(n9191) );
  NAND2X0_RVT U8876 ( .A1(n5272), .A2(n7009), .Y(n7047) );
  NAND3X0_RVT U8877 ( .A1(n9232), .A2(n6432), .A3(n9233), .Y(n8673) );
  NAND2X0_RVT U8878 ( .A1(n8881), .A2(n5265), .Y(n9233) );
  NAND3X0_RVT U8879 ( .A1(n6739), .A2(n5271), .A3(n5272), .Y(n8507) );
  INVX0_RVT U8880 ( .A(n9234), .Y(n5272) );
  NAND3X0_RVT U8881 ( .A1(n4905), .A2(n4910), .A3(n8560), .Y(n6432) );
  AND2X1_RVT U8882 ( .A1(n792), .A2(n789), .Y(n8560) );
  NAND3X0_RVT U8883 ( .A1(n7009), .A2(n5271), .A3(n8510), .Y(n9232) );
  INVX0_RVT U8884 ( .A(n5270), .Y(n8510) );
  NAND2X0_RVT U8885 ( .A1(n5301), .A2(n5280), .Y(n5271) );
  NAND3X0_RVT U8886 ( .A1(n731), .A2(n4913), .A3(n732), .Y(n5280) );
  AND2X1_RVT U8887 ( .A1(n5265), .A2(n6739), .Y(n7009) );
  NAND2X0_RVT U8888 ( .A1(n9235), .A2(n9236), .Y(n6739) );
  NAND2X0_RVT U8889 ( .A1(n8491), .A2(n9237), .Y(n9236) );
  INVX0_RVT U8890 ( .A(n6476), .Y(n8491) );
  NAND2X0_RVT U8891 ( .A1(n9238), .A2(n9239), .Y(n9235) );
  NAND2X0_RVT U8892 ( .A1(n9240), .A2(n9241), .Y(n9239) );
  NAND2X0_RVT U8893 ( .A1(n9242), .A2(n6476), .Y(n9241) );
  NAND2X0_RVT U8894 ( .A1(n9243), .A2(n9244), .Y(n9240) );
  NAND3X0_RVT U8895 ( .A1(n9245), .A2(n9246), .A3(n9247), .Y(n9244) );
  OR2X1_RVT U8896 ( .A1(n9248), .A2(n9249), .Y(n9247) );
  NAND2X0_RVT U8897 ( .A1(n9250), .A2(n6476), .Y(n9246) );
  NAND4X0_RVT U8898 ( .A1(n7912), .A2(n6756), .A3(n9251), .A4(n6476), .Y(n9245) );
  NAND2X0_RVT U8899 ( .A1(n9249), .A2(n9248), .Y(n9243) );
  NAND2X0_RVT U8900 ( .A1(n6738), .A2(n6743), .Y(n9248) );
  INVX0_RVT U8901 ( .A(n8517), .Y(n6738) );
  NAND2X0_RVT U8902 ( .A1(n9121), .A2(n6727), .Y(n8517) );
  NAND2X0_RVT U8903 ( .A1(n9252), .A2(n6476), .Y(n9249) );
  INVX0_RVT U8904 ( .A(n9237), .Y(n9238) );
  NAND2X0_RVT U8905 ( .A1(n9253), .A2(n9254), .Y(n9237) );
  NAND2X0_RVT U8906 ( .A1(n8515), .A2(n8182), .Y(n9254) );
  NAND4X0_RVT U8907 ( .A1(n9255), .A2(n9256), .A3(n9257), .A4(n9258), .Y(n8182) );
  NAND2X0_RVT U8908 ( .A1(n7842), .A2(n9259), .Y(n9258) );
  NAND4X0_RVT U8909 ( .A1(n9260), .A2(n9261), .A3(n9262), .A4(n9263), .Y(n9259) );
  NAND2X0_RVT U8910 ( .A1(n7694), .A2(n5167), .Y(n9263) );
  NAND2X0_RVT U8911 ( .A1(n7678), .A2(n5043), .Y(n9262) );
  NAND2X0_RVT U8912 ( .A1(n7766), .A2(n5044), .Y(n9261) );
  NAND2X0_RVT U8913 ( .A1(n8501), .A2(n5045), .Y(n9260) );
  NAND2X0_RVT U8914 ( .A1(n7853), .A2(n9129), .Y(n9257) );
  NAND4X0_RVT U8915 ( .A1(n9264), .A2(n9265), .A3(n9266), .A4(n9267), .Y(n9129) );
  NAND2X0_RVT U8916 ( .A1(n7694), .A2(n5168), .Y(n9267) );
  NAND2X0_RVT U8917 ( .A1(n7678), .A2(n5046), .Y(n9266) );
  NAND2X0_RVT U8918 ( .A1(n7766), .A2(n5047), .Y(n9265) );
  NAND2X0_RVT U8919 ( .A1(n8501), .A2(n5048), .Y(n9264) );
  NAND2X0_RVT U8920 ( .A1(n7848), .A2(n7750), .Y(n9256) );
  NAND4X0_RVT U8921 ( .A1(n9268), .A2(n9269), .A3(n9270), .A4(n9271), .Y(n7750) );
  NAND2X0_RVT U8922 ( .A1(n7694), .A2(n5169), .Y(n9271) );
  NAND2X0_RVT U8923 ( .A1(n7678), .A2(n5170), .Y(n9270) );
  NAND2X0_RVT U8924 ( .A1(n7766), .A2(n5171), .Y(n9269) );
  NAND2X0_RVT U8925 ( .A1(n8501), .A2(n5049), .Y(n9268) );
  NAND2X0_RVT U8926 ( .A1(n7852), .A2(n7753), .Y(n9255) );
  NAND4X0_RVT U8927 ( .A1(n9272), .A2(n9273), .A3(n9274), .A4(n9275), .Y(n7753) );
  NAND2X0_RVT U8928 ( .A1(n7694), .A2(n5172), .Y(n9275) );
  NAND2X0_RVT U8929 ( .A1(n7678), .A2(n5050), .Y(n9274) );
  NAND2X0_RVT U8930 ( .A1(n7766), .A2(n5051), .Y(n9273) );
  NAND2X0_RVT U8931 ( .A1(n8501), .A2(n5194), .Y(n9272) );
  AND2X1_RVT U8932 ( .A1(n4906), .A2(n4926), .Y(n8501) );
  INVX0_RVT U8933 ( .A(n6434), .Y(n8515) );
  NAND2X0_RVT U8934 ( .A1(n9276), .A2(n9277), .Y(n6434) );
  NAND2X0_RVT U8935 ( .A1(n6736), .A2(n9278), .Y(n9277) );
  NAND2X0_RVT U8936 ( .A1(n9242), .A2(n6736), .Y(n9281) );
  AND3X1_RVT U8937 ( .A1(n9282), .A2(n4930), .A3(n936), .Y(n9242) );
  NAND2X0_RVT U8938 ( .A1(n6736), .A2(n9252), .Y(n9280) );
  XNOR3X1_RVT U8939 ( .A1(n4907), .A2(n937), .A3(n9283), .Y(n9252) );
  NAND3X0_RVT U8940 ( .A1(n9250), .A2(n9251), .A3(n6736), .Y(n9279) );
  NOR2X0_RVT U8941 ( .A1(n6407), .A2(n6453), .Y(n6736) );
  NAND2X0_RVT U8942 ( .A1(n9284), .A2(n9285), .Y(n6453) );
  NAND2X0_RVT U8943 ( .A1(n9286), .A2(n9287), .Y(n9251) );
  NAND2X0_RVT U8944 ( .A1(n939), .A2(n4928), .Y(n9287) );
  XNOR3X1_RVT U8945 ( .A1(n4909), .A2(n938), .A3(n9288), .Y(n9250) );
  INVX0_RVT U8946 ( .A(n5340), .Y(n6306) );
  NAND3X0_RVT U8947 ( .A1(n6760), .A2(n4925), .A3(n792), .Y(n5340) );
  AND2X1_RVT U8948 ( .A1(n790), .A2(n791), .Y(n6760) );
  NAND2X0_RVT U8949 ( .A1(n9278), .A2(n6476), .Y(n9253) );
  NAND3X0_RVT U8950 ( .A1(n6743), .A2(n6727), .A3(n6509), .Y(n6476) );
  AND3X1_RVT U8951 ( .A1(n6756), .A2(n9121), .A3(n7912), .Y(n6509) );
  INVX0_RVT U8952 ( .A(n7279), .Y(n7912) );
  NAND2X0_RVT U8953 ( .A1(n7010), .A2(n5270), .Y(n7279) );
  NAND2X0_RVT U8954 ( .A1(n9289), .A2(n6330), .Y(n5270) );
  NAND2X0_RVT U8955 ( .A1(n8512), .A2(n9289), .Y(n7010) );
  AND4X1_RVT U8956 ( .A1(n8514), .A2(n9230), .A3(n9285), .A4(n6339), .Y(n9289)
         );
  INVX0_RVT U8957 ( .A(n6348), .Y(n9230) );
  NAND3X0_RVT U8958 ( .A1(n8514), .A2(n9290), .A3(n9291), .Y(n9121) );
  INVX0_RVT U8959 ( .A(n6321), .Y(n8514) );
  AND2X1_RVT U8960 ( .A1(n9234), .A2(n8511), .Y(n6756) );
  NAND2X0_RVT U8961 ( .A1(n9292), .A2(n9284), .Y(n8511) );
  NAND3X0_RVT U8962 ( .A1(n9290), .A2(n6321), .A3(n9292), .Y(n9234) );
  AND3X1_RVT U8963 ( .A1(n9227), .A2(n9293), .A3(n9229), .Y(n9292) );
  INVX0_RVT U8964 ( .A(n6370), .Y(n9229) );
  NAND2X0_RVT U8965 ( .A1(n9291), .A2(n9284), .Y(n6727) );
  AND4X1_RVT U8966 ( .A1(n9231), .A2(n6321), .A3(n6348), .A4(n6330), .Y(n9284)
         );
  AND3X1_RVT U8967 ( .A1(n6370), .A2(n6358), .A3(n9293), .Y(n9291) );
  NOR2X0_RVT U8968 ( .A1(n6387), .A2(n9228), .Y(n9293) );
  INVX0_RVT U8969 ( .A(n6307), .Y(n9228) );
  NAND3X0_RVT U8970 ( .A1(n9285), .A2(n6321), .A3(n9290), .Y(n6743) );
  AND3X1_RVT U8971 ( .A1(n9231), .A2(n6348), .A3(n8512), .Y(n9290) );
  INVX0_RVT U8972 ( .A(n6330), .Y(n8512) );
  NAND2X0_RVT U8973 ( .A1(n9294), .A2(n9295), .Y(n6330) );
  OR3X1_RVT U8974 ( .A1(n9296), .A2(n9297), .A3(n936), .Y(n9295) );
  NAND4X0_RVT U8975 ( .A1(n9298), .A2(n9299), .A3(n9300), .A4(n9301), .Y(n9297) );
  NAND2X0_RVT U8976 ( .A1(n862), .A2(n9302), .Y(n9301) );
  NAND2X0_RVT U8977 ( .A1(n854), .A2(n9303), .Y(n9300) );
  NAND2X0_RVT U8978 ( .A1(n846), .A2(n9304), .Y(n9299) );
  NAND2X0_RVT U8979 ( .A1(n830), .A2(n9305), .Y(n9298) );
  NAND4X0_RVT U8980 ( .A1(n9306), .A2(n9307), .A3(n9308), .A4(n9309), .Y(n9296) );
  NAND2X0_RVT U8981 ( .A1(n822), .A2(n9310), .Y(n9309) );
  NAND2X0_RVT U8982 ( .A1(n838), .A2(n9311), .Y(n9308) );
  NAND2X0_RVT U8983 ( .A1(n813), .A2(n9312), .Y(n9307) );
  NAND2X0_RVT U8984 ( .A1(n870), .A2(n9313), .Y(n9306) );
  OR3X1_RVT U8985 ( .A1(n9314), .A2(n9315), .A3(n4906), .Y(n9294) );
  NAND4X0_RVT U8986 ( .A1(n9316), .A2(n9317), .A3(n9318), .A4(n9319), .Y(n9315) );
  NAND2X0_RVT U8987 ( .A1(n926), .A2(n9302), .Y(n9319) );
  NAND2X0_RVT U8988 ( .A1(n918), .A2(n9303), .Y(n9318) );
  NAND2X0_RVT U8989 ( .A1(n910), .A2(n9304), .Y(n9317) );
  NAND2X0_RVT U8990 ( .A1(n894), .A2(n9305), .Y(n9316) );
  NAND4X0_RVT U8991 ( .A1(n9320), .A2(n9321), .A3(n9322), .A4(n9323), .Y(n9314) );
  NAND2X0_RVT U8992 ( .A1(n886), .A2(n9310), .Y(n9323) );
  NAND2X0_RVT U8993 ( .A1(n902), .A2(n9311), .Y(n9322) );
  NAND2X0_RVT U8994 ( .A1(n878), .A2(n9312), .Y(n9321) );
  NAND2X0_RVT U8995 ( .A1(n934), .A2(n9313), .Y(n9320) );
  NAND2X0_RVT U8996 ( .A1(n9324), .A2(n9325), .Y(n6348) );
  OR3X1_RVT U8997 ( .A1(n9326), .A2(n9327), .A3(n936), .Y(n9325) );
  NAND4X0_RVT U8998 ( .A1(n9328), .A2(n9329), .A3(n9330), .A4(n9331), .Y(n9327) );
  NAND2X0_RVT U8999 ( .A1(n860), .A2(n9302), .Y(n9331) );
  NAND2X0_RVT U9000 ( .A1(n852), .A2(n9303), .Y(n9330) );
  NAND2X0_RVT U9001 ( .A1(n844), .A2(n9304), .Y(n9329) );
  NAND2X0_RVT U9002 ( .A1(n828), .A2(n9305), .Y(n9328) );
  NAND4X0_RVT U9003 ( .A1(n9332), .A2(n9333), .A3(n9334), .A4(n9335), .Y(n9326) );
  NAND2X0_RVT U9004 ( .A1(n820), .A2(n9310), .Y(n9335) );
  NAND2X0_RVT U9005 ( .A1(n836), .A2(n9311), .Y(n9334) );
  NAND2X0_RVT U9006 ( .A1(n809), .A2(n9312), .Y(n9333) );
  NAND2X0_RVT U9007 ( .A1(n868), .A2(n9313), .Y(n9332) );
  OR3X1_RVT U9008 ( .A1(n9336), .A2(n9337), .A3(n4906), .Y(n9324) );
  NAND4X0_RVT U9009 ( .A1(n9338), .A2(n9339), .A3(n9340), .A4(n9341), .Y(n9337) );
  NAND2X0_RVT U9010 ( .A1(n924), .A2(n9302), .Y(n9341) );
  NAND2X0_RVT U9011 ( .A1(n916), .A2(n9303), .Y(n9340) );
  NAND2X0_RVT U9012 ( .A1(n908), .A2(n9304), .Y(n9339) );
  NAND2X0_RVT U9013 ( .A1(n892), .A2(n9305), .Y(n9338) );
  NAND4X0_RVT U9014 ( .A1(n9342), .A2(n9343), .A3(n9344), .A4(n9345), .Y(n9336) );
  NAND2X0_RVT U9015 ( .A1(n884), .A2(n9310), .Y(n9345) );
  NAND2X0_RVT U9016 ( .A1(n900), .A2(n9311), .Y(n9344) );
  NAND2X0_RVT U9017 ( .A1(n876), .A2(n9312), .Y(n9343) );
  NAND2X0_RVT U9018 ( .A1(n932), .A2(n9313), .Y(n9342) );
  INVX0_RVT U9019 ( .A(n6339), .Y(n9231) );
  NAND2X0_RVT U9020 ( .A1(n9346), .A2(n9347), .Y(n6339) );
  OR3X1_RVT U9021 ( .A1(n9348), .A2(n9349), .A3(n936), .Y(n9347) );
  NAND4X0_RVT U9022 ( .A1(n9350), .A2(n9351), .A3(n9352), .A4(n9353), .Y(n9349) );
  NAND2X0_RVT U9023 ( .A1(n861), .A2(n9302), .Y(n9353) );
  NAND2X0_RVT U9024 ( .A1(n853), .A2(n9303), .Y(n9352) );
  NAND2X0_RVT U9025 ( .A1(n845), .A2(n9304), .Y(n9351) );
  NAND2X0_RVT U9026 ( .A1(n829), .A2(n9305), .Y(n9350) );
  NAND4X0_RVT U9027 ( .A1(n9354), .A2(n9355), .A3(n9356), .A4(n9357), .Y(n9348) );
  NAND2X0_RVT U9028 ( .A1(n821), .A2(n9310), .Y(n9357) );
  NAND2X0_RVT U9029 ( .A1(n837), .A2(n9311), .Y(n9356) );
  NAND2X0_RVT U9030 ( .A1(n811), .A2(n9312), .Y(n9355) );
  NAND2X0_RVT U9031 ( .A1(n869), .A2(n9313), .Y(n9354) );
  OR3X1_RVT U9032 ( .A1(n9358), .A2(n9359), .A3(n4906), .Y(n9346) );
  NAND4X0_RVT U9033 ( .A1(n9360), .A2(n9361), .A3(n9362), .A4(n9363), .Y(n9359) );
  NAND2X0_RVT U9034 ( .A1(n925), .A2(n9302), .Y(n9363) );
  NAND2X0_RVT U9035 ( .A1(n917), .A2(n9303), .Y(n9362) );
  NAND2X0_RVT U9036 ( .A1(n909), .A2(n9304), .Y(n9361) );
  NAND2X0_RVT U9037 ( .A1(n893), .A2(n9305), .Y(n9360) );
  NAND4X0_RVT U9038 ( .A1(n9364), .A2(n9365), .A3(n9366), .A4(n9367), .Y(n9358) );
  NAND2X0_RVT U9039 ( .A1(n885), .A2(n9310), .Y(n9367) );
  NAND2X0_RVT U9040 ( .A1(n901), .A2(n9311), .Y(n9366) );
  NAND2X0_RVT U9041 ( .A1(n877), .A2(n9312), .Y(n9365) );
  NAND2X0_RVT U9042 ( .A1(n933), .A2(n9313), .Y(n9364) );
  NAND2X0_RVT U9043 ( .A1(n9368), .A2(n9369), .Y(n6321) );
  OR3X1_RVT U9044 ( .A1(n9370), .A2(n9371), .A3(n936), .Y(n9369) );
  NAND4X0_RVT U9045 ( .A1(n9372), .A2(n9373), .A3(n9374), .A4(n9375), .Y(n9371) );
  NAND2X0_RVT U9046 ( .A1(n863), .A2(n9302), .Y(n9375) );
  NAND2X0_RVT U9047 ( .A1(n855), .A2(n9303), .Y(n9374) );
  NAND2X0_RVT U9048 ( .A1(n847), .A2(n9304), .Y(n9373) );
  NAND2X0_RVT U9049 ( .A1(n831), .A2(n9305), .Y(n9372) );
  NAND4X0_RVT U9050 ( .A1(n9376), .A2(n9377), .A3(n9378), .A4(n9379), .Y(n9370) );
  NAND2X0_RVT U9051 ( .A1(n823), .A2(n9310), .Y(n9379) );
  NAND2X0_RVT U9052 ( .A1(n839), .A2(n9311), .Y(n9378) );
  NAND2X0_RVT U9053 ( .A1(n815), .A2(n9312), .Y(n9377) );
  NAND2X0_RVT U9054 ( .A1(n871), .A2(n9313), .Y(n9376) );
  OR3X1_RVT U9055 ( .A1(n9380), .A2(n9381), .A3(n4906), .Y(n9368) );
  NAND4X0_RVT U9056 ( .A1(n9382), .A2(n9383), .A3(n9384), .A4(n9385), .Y(n9381) );
  NAND2X0_RVT U9057 ( .A1(n927), .A2(n9302), .Y(n9385) );
  NAND2X0_RVT U9058 ( .A1(n919), .A2(n9303), .Y(n9384) );
  NAND2X0_RVT U9059 ( .A1(n911), .A2(n9304), .Y(n9383) );
  NAND2X0_RVT U9060 ( .A1(n895), .A2(n9305), .Y(n9382) );
  NAND4X0_RVT U9061 ( .A1(n9386), .A2(n9387), .A3(n9388), .A4(n9389), .Y(n9380) );
  NAND2X0_RVT U9062 ( .A1(n887), .A2(n9310), .Y(n9389) );
  NAND2X0_RVT U9063 ( .A1(n903), .A2(n9311), .Y(n9388) );
  NAND2X0_RVT U9064 ( .A1(n879), .A2(n9312), .Y(n9387) );
  NAND2X0_RVT U9065 ( .A1(n935), .A2(n9313), .Y(n9386) );
  AND4X1_RVT U9066 ( .A1(n9227), .A2(n6370), .A3(n6307), .A4(n6387), .Y(n9285)
         );
  NAND2X0_RVT U9067 ( .A1(n9390), .A2(n9391), .Y(n6387) );
  OR3X1_RVT U9068 ( .A1(n9392), .A2(n9393), .A3(n936), .Y(n9391) );
  NAND4X0_RVT U9069 ( .A1(n9394), .A2(n9395), .A3(n9396), .A4(n9397), .Y(n9393) );
  NAND2X0_RVT U9070 ( .A1(n857), .A2(n9302), .Y(n9397) );
  NAND2X0_RVT U9071 ( .A1(n849), .A2(n9303), .Y(n9396) );
  NAND2X0_RVT U9072 ( .A1(n841), .A2(n9304), .Y(n9395) );
  NAND2X0_RVT U9073 ( .A1(n825), .A2(n9305), .Y(n9394) );
  NAND4X0_RVT U9074 ( .A1(n9398), .A2(n9399), .A3(n9400), .A4(n9401), .Y(n9392) );
  NAND2X0_RVT U9075 ( .A1(n817), .A2(n9310), .Y(n9401) );
  NAND2X0_RVT U9076 ( .A1(n833), .A2(n9311), .Y(n9400) );
  NAND2X0_RVT U9077 ( .A1(n803), .A2(n9312), .Y(n9399) );
  NAND2X0_RVT U9078 ( .A1(n865), .A2(n9313), .Y(n9398) );
  OR3X1_RVT U9079 ( .A1(n9402), .A2(n9403), .A3(n4906), .Y(n9390) );
  NAND4X0_RVT U9080 ( .A1(n9404), .A2(n9405), .A3(n9406), .A4(n9407), .Y(n9403) );
  NAND2X0_RVT U9081 ( .A1(n921), .A2(n9302), .Y(n9407) );
  NAND2X0_RVT U9082 ( .A1(n913), .A2(n9303), .Y(n9406) );
  NAND2X0_RVT U9083 ( .A1(n905), .A2(n9304), .Y(n9405) );
  NAND2X0_RVT U9084 ( .A1(n889), .A2(n9305), .Y(n9404) );
  NAND4X0_RVT U9085 ( .A1(n9408), .A2(n9409), .A3(n9410), .A4(n9411), .Y(n9402) );
  NAND2X0_RVT U9086 ( .A1(n881), .A2(n9310), .Y(n9411) );
  NAND2X0_RVT U9087 ( .A1(n897), .A2(n9311), .Y(n9410) );
  NAND2X0_RVT U9088 ( .A1(n873), .A2(n9312), .Y(n9409) );
  NAND2X0_RVT U9089 ( .A1(n929), .A2(n9313), .Y(n9408) );
  NAND2X0_RVT U9090 ( .A1(n9412), .A2(n9413), .Y(n6307) );
  OR3X1_RVT U9091 ( .A1(n9414), .A2(n9415), .A3(n936), .Y(n9413) );
  NAND4X0_RVT U9092 ( .A1(n9416), .A2(n9417), .A3(n9418), .A4(n9419), .Y(n9415) );
  NAND2X0_RVT U9093 ( .A1(n856), .A2(n9302), .Y(n9419) );
  NAND2X0_RVT U9094 ( .A1(n848), .A2(n9303), .Y(n9418) );
  NAND2X0_RVT U9095 ( .A1(n840), .A2(n9304), .Y(n9417) );
  NAND2X0_RVT U9096 ( .A1(n824), .A2(n9305), .Y(n9416) );
  NAND4X0_RVT U9097 ( .A1(n9420), .A2(n9421), .A3(n9422), .A4(n9423), .Y(n9414) );
  NAND2X0_RVT U9098 ( .A1(n816), .A2(n9310), .Y(n9423) );
  NAND2X0_RVT U9099 ( .A1(n832), .A2(n9311), .Y(n9422) );
  NAND2X0_RVT U9100 ( .A1(n801), .A2(n9312), .Y(n9421) );
  NAND2X0_RVT U9101 ( .A1(n864), .A2(n9313), .Y(n9420) );
  OR3X1_RVT U9102 ( .A1(n9424), .A2(n9425), .A3(n4906), .Y(n9412) );
  NAND4X0_RVT U9103 ( .A1(n9426), .A2(n9427), .A3(n9428), .A4(n9429), .Y(n9425) );
  NAND2X0_RVT U9104 ( .A1(n920), .A2(n9302), .Y(n9429) );
  NAND2X0_RVT U9105 ( .A1(n912), .A2(n9303), .Y(n9428) );
  NAND2X0_RVT U9106 ( .A1(n904), .A2(n9304), .Y(n9427) );
  NAND2X0_RVT U9107 ( .A1(n888), .A2(n9305), .Y(n9426) );
  NAND4X0_RVT U9108 ( .A1(n9430), .A2(n9431), .A3(n9432), .A4(n9433), .Y(n9424) );
  NAND2X0_RVT U9109 ( .A1(n880), .A2(n9310), .Y(n9433) );
  NAND2X0_RVT U9110 ( .A1(n896), .A2(n9311), .Y(n9432) );
  NAND2X0_RVT U9111 ( .A1(n872), .A2(n9312), .Y(n9431) );
  NAND2X0_RVT U9112 ( .A1(n928), .A2(n9313), .Y(n9430) );
  NAND2X0_RVT U9113 ( .A1(n9434), .A2(n9435), .Y(n6370) );
  OR3X1_RVT U9114 ( .A1(n9436), .A2(n9437), .A3(n936), .Y(n9435) );
  NAND4X0_RVT U9115 ( .A1(n9438), .A2(n9439), .A3(n9440), .A4(n9441), .Y(n9437) );
  NAND2X0_RVT U9116 ( .A1(n858), .A2(n9302), .Y(n9441) );
  NAND2X0_RVT U9117 ( .A1(n850), .A2(n9303), .Y(n9440) );
  NAND2X0_RVT U9118 ( .A1(n842), .A2(n9304), .Y(n9439) );
  NAND2X0_RVT U9119 ( .A1(n826), .A2(n9305), .Y(n9438) );
  NAND4X0_RVT U9120 ( .A1(n9442), .A2(n9443), .A3(n9444), .A4(n9445), .Y(n9436) );
  NAND2X0_RVT U9121 ( .A1(n818), .A2(n9310), .Y(n9445) );
  NAND2X0_RVT U9122 ( .A1(n834), .A2(n9311), .Y(n9444) );
  NAND2X0_RVT U9123 ( .A1(n805), .A2(n9312), .Y(n9443) );
  NAND2X0_RVT U9124 ( .A1(n866), .A2(n9313), .Y(n9442) );
  OR3X1_RVT U9125 ( .A1(n9446), .A2(n9447), .A3(n4906), .Y(n9434) );
  NAND4X0_RVT U9126 ( .A1(n9448), .A2(n9449), .A3(n9450), .A4(n9451), .Y(n9447) );
  NAND2X0_RVT U9127 ( .A1(n922), .A2(n9302), .Y(n9451) );
  NAND2X0_RVT U9128 ( .A1(n914), .A2(n9303), .Y(n9450) );
  NAND2X0_RVT U9129 ( .A1(n906), .A2(n9304), .Y(n9449) );
  NAND2X0_RVT U9130 ( .A1(n890), .A2(n9305), .Y(n9448) );
  NAND4X0_RVT U9131 ( .A1(n9452), .A2(n9453), .A3(n9454), .A4(n9455), .Y(n9446) );
  NAND2X0_RVT U9132 ( .A1(n882), .A2(n9310), .Y(n9455) );
  NAND2X0_RVT U9133 ( .A1(n898), .A2(n9311), .Y(n9454) );
  NAND2X0_RVT U9134 ( .A1(n874), .A2(n9312), .Y(n9453) );
  NAND2X0_RVT U9135 ( .A1(n930), .A2(n9313), .Y(n9452) );
  INVX0_RVT U9136 ( .A(n6358), .Y(n9227) );
  NAND2X0_RVT U9137 ( .A1(n9456), .A2(n9457), .Y(n6358) );
  OR3X1_RVT U9138 ( .A1(n9458), .A2(n9459), .A3(n936), .Y(n9457) );
  NAND4X0_RVT U9139 ( .A1(n9460), .A2(n9461), .A3(n9462), .A4(n9463), .Y(n9459) );
  NAND2X0_RVT U9140 ( .A1(n859), .A2(n9302), .Y(n9463) );
  NAND2X0_RVT U9141 ( .A1(n851), .A2(n9303), .Y(n9462) );
  NAND2X0_RVT U9142 ( .A1(n843), .A2(n9304), .Y(n9461) );
  NAND2X0_RVT U9143 ( .A1(n827), .A2(n9305), .Y(n9460) );
  NAND4X0_RVT U9144 ( .A1(n9464), .A2(n9465), .A3(n9466), .A4(n9467), .Y(n9458) );
  NAND2X0_RVT U9145 ( .A1(n819), .A2(n9310), .Y(n9467) );
  NAND2X0_RVT U9146 ( .A1(n835), .A2(n9311), .Y(n9466) );
  NAND2X0_RVT U9147 ( .A1(n807), .A2(n9312), .Y(n9465) );
  NAND2X0_RVT U9148 ( .A1(n867), .A2(n9313), .Y(n9464) );
  OR3X1_RVT U9149 ( .A1(n9468), .A2(n9469), .A3(n4906), .Y(n9456) );
  NAND4X0_RVT U9150 ( .A1(n9470), .A2(n9471), .A3(n9472), .A4(n9473), .Y(n9469) );
  NAND2X0_RVT U9151 ( .A1(n923), .A2(n9302), .Y(n9473) );
  AND2X1_RVT U9152 ( .A1(n7853), .A2(n937), .Y(n9302) );
  NAND2X0_RVT U9153 ( .A1(n915), .A2(n9303), .Y(n9472) );
  AND2X1_RVT U9154 ( .A1(n937), .A2(n7852), .Y(n9303) );
  NAND2X0_RVT U9155 ( .A1(n907), .A2(n9304), .Y(n9471) );
  AND2X1_RVT U9156 ( .A1(n937), .A2(n7848), .Y(n9304) );
  NAND2X0_RVT U9157 ( .A1(n891), .A2(n9305), .Y(n9470) );
  AND2X1_RVT U9158 ( .A1(n7853), .A2(n4926), .Y(n9305) );
  NAND4X0_RVT U9159 ( .A1(n9474), .A2(n9475), .A3(n9476), .A4(n9477), .Y(n9468) );
  NAND2X0_RVT U9160 ( .A1(n883), .A2(n9310), .Y(n9477) );
  AND2X1_RVT U9161 ( .A1(n7852), .A2(n4926), .Y(n9310) );
  NAND2X0_RVT U9162 ( .A1(n899), .A2(n9311), .Y(n9476) );
  AND2X1_RVT U9163 ( .A1(n7842), .A2(n4926), .Y(n9311) );
  NAND2X0_RVT U9164 ( .A1(n875), .A2(n9312), .Y(n9475) );
  AND2X1_RVT U9165 ( .A1(n7848), .A2(n4926), .Y(n9312) );
  NAND2X0_RVT U9166 ( .A1(n931), .A2(n9313), .Y(n9474) );
  AND2X1_RVT U9167 ( .A1(n937), .A2(n7842), .Y(n9313) );
  NAND2X0_RVT U9168 ( .A1(n9479), .A2(n9480), .Y(n9478) );
  NAND2X0_RVT U9169 ( .A1(n9481), .A2(n4930), .Y(n9480) );
  OR2X1_RVT U9170 ( .A1(n9282), .A2(n936), .Y(n9481) );
  NAND2X0_RVT U9171 ( .A1(n936), .A2(n9282), .Y(n9479) );
  NAND2X0_RVT U9172 ( .A1(n9482), .A2(n9483), .Y(n9282) );
  NAND2X0_RVT U9173 ( .A1(n9484), .A2(n4907), .Y(n9483) );
  NAND2X0_RVT U9174 ( .A1(n9283), .A2(n4926), .Y(n9484) );
  INVX0_RVT U9175 ( .A(n9485), .Y(n9283) );
  NAND2X0_RVT U9176 ( .A1(n937), .A2(n9485), .Y(n9482) );
  NAND2X0_RVT U9177 ( .A1(n9486), .A2(n9487), .Y(n9485) );
  NAND2X0_RVT U9178 ( .A1(n9488), .A2(n4909), .Y(n9487) );
  NAND2X0_RVT U9179 ( .A1(n9288), .A2(n4927), .Y(n9488) );
  INVX0_RVT U9180 ( .A(n9286), .Y(n9288) );
  NAND2X0_RVT U9181 ( .A1(n938), .A2(n9286), .Y(n9486) );
  NAND2X0_RVT U9182 ( .A1(n975), .A2(n4908), .Y(n9286) );
  NAND3X0_RVT U9183 ( .A1(n6534), .A2(n4905), .A3(n791), .Y(n6407) );
  AND2X1_RVT U9184 ( .A1(n789), .A2(n4969), .Y(n6534) );
  NAND3X0_RVT U9185 ( .A1(n9489), .A2(n9490), .A3(n9491), .Y(n4495) );
  NAND2X0_RVT U9186 ( .A1(n9492), .A2(n5190), .Y(n9491) );
  NAND2X0_RVT U9187 ( .A1(n9514), .A2(n5053), .Y(n9489) );
  NAND2X0_RVT U9188 ( .A1(n9493), .A2(n9494), .Y(n4494) );
  NAND2X0_RVT U9189 ( .A1(n5276), .A2(BE_n[3]), .Y(n9494) );
  NAND2X0_RVT U9190 ( .A1(n6751), .A2(n5190), .Y(n9493) );
  NAND3X0_RVT U9191 ( .A1(n9495), .A2(n9496), .A3(n9497), .Y(n4493) );
  NAND2X0_RVT U9192 ( .A1(n9492), .A2(n5191), .Y(n9497) );
  NAND3X0_RVT U9193 ( .A1(n9498), .A2(n5053), .A3(n9514), .Y(n9496) );
  NAND2X0_RVT U9194 ( .A1(rEIP[0]), .A2(n4914), .Y(n9498) );
  NAND2X0_RVT U9195 ( .A1(n9499), .A2(rEIP[0]), .Y(n9495) );
  INVX0_RVT U9196 ( .A(n9500), .Y(n9499) );
  NAND2X0_RVT U9197 ( .A1(n9501), .A2(n9502), .Y(n4492) );
  NAND2X0_RVT U9198 ( .A1(n5276), .A2(BE_n[2]), .Y(n9502) );
  NAND2X0_RVT U9199 ( .A1(n6751), .A2(n5191), .Y(n9501) );
  NAND3X0_RVT U9200 ( .A1(n9500), .A2(n9490), .A3(n9503), .Y(n4491) );
  NAND2X0_RVT U9201 ( .A1(n9492), .A2(n5192), .Y(n9503) );
  OR3X1_RVT U9202 ( .A1(n4914), .A2(rEIP[0]), .A3(n4968), .Y(n9490) );
  NAND2X0_RVT U9203 ( .A1(n9504), .A2(n9505), .Y(n4490) );
  NAND2X0_RVT U9204 ( .A1(n5276), .A2(BE_n[1]), .Y(n9505) );
  NAND2X0_RVT U9205 ( .A1(n6751), .A2(n5192), .Y(n9504) );
  NAND3X0_RVT U9206 ( .A1(n9506), .A2(n9507), .A3(n9500), .Y(n4489) );
  NAND2X0_RVT U9207 ( .A1(rEIP[1]), .A2(n9508), .Y(n9500) );
  NAND2X0_RVT U9208 ( .A1(n9492), .A2(n5193), .Y(n9507) );
  INVX0_RVT U9209 ( .A(n9508), .Y(n9492) );
  NAND2X0_RVT U9210 ( .A1(rEIP[0]), .A2(n9508), .Y(n9506) );
  NAND2X0_RVT U9211 ( .A1(n4914), .A2(n4968), .Y(n9508) );
  NAND2X0_RVT U9212 ( .A1(n9509), .A2(n9510), .Y(n4488) );
  NAND2X0_RVT U9213 ( .A1(n5276), .A2(BE_n[0]), .Y(n9510) );
  NAND2X0_RVT U9214 ( .A1(n6751), .A2(n5193), .Y(n9509) );
  NAND2X0_RVT U9215 ( .A1(n5301), .A2(n5279), .Y(n6751) );
  NAND3X0_RVT U9216 ( .A1(n4913), .A2(n4962), .A3(n732), .Y(n5279) );
  NAND2X0_RVT U9217 ( .A1(n5296), .A2(n732), .Y(n5301) );
  INVX0_RVT U9218 ( .A(n5278), .Y(n5296) );
  NAND2X0_RVT U9219 ( .A1(n730), .A2(n4962), .Y(n5278) );
  //new;
endmodule