
module c432 ( N1, N4, N8, N11, N14, N17, N21, N24, N27, N30, N34, N37, N40, 
        N43, N47, N50, N53, N56, N60, N63, N66, N69, N73, N76, N79, N82, N86, 
        N89, N92, N95, N99, N102, N105, N108, N112, N115, N223, N329, N370, 
        N421, N430, N431, N432 );
  input N1, N4, N8, N11, N14, N17, N21, N24, N27, N30, N34, N37, N40, N43, N47, N50, N53, N56, N60, N63, N66, N69, N73, N76, N79, N82, N86, N89, N92, N95, N99, N102, N105, N108, N112, N115;
  output N223, N329, N370, N421, N430, N431, N432;
  wire   n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257;
n60001, n60002, n60003, n60004, n60005, n60006, n60007, n60008, n60009, n60010;
//add;

//gate;
NAND2X0_RVT U134 ( .A1(n133), .A2(n134), .Y(N432) );
  AND2X0_RVT U135 ( .A1(n135), .A2(n136), .Y(n60001) );
  NAND3X0_RVT U136 ( .A1(n137), .A2(n138), .A3(n139), .Y(n135) );
  NAND2X0_RVT U137 ( .A1(n140), .A2(n141), .Y(n139) );
  INVX0_RVT U138 ( .A(n142), .Y(n140) );
  NAND4X0_RVT U139 ( .A1(n143), .A2(n144), .A3(n145), .A4(n146), .Y(n137) );
  NAND2X0_RVT U140 ( .A1(N99), .A2(N329), .Y(n144) );
  NAND2X0_RVT U141 ( .A1(N105), .A2(N370), .Y(n60007) );
  NAND3X0_RVT U142 ( .A1(n133), .A2(n136), .A3(n147), .Y(N431) );
  NAND3X0_RVT U143 ( .A1(n138), .A2(n141), .A3(n148), .Y(n147) );
  AND2X1_RVT U144 ( .A1(n149), .A2(n150), .Y(N421) );
  OR4X1_RVT U145 ( .A1(n145), .A2(n148), .A3(N430), .A4(N108), .Y(n150) );
  NAND4X0_RVT U146 ( .A1(n138), .A2(n141), .A3(n133), .A4(n136), .Y(N430) );
  NAND3X0_RVT U147 ( .A1(n151), .A2(n152), .A3(n153), .Y(n136) );
  NAND2X0_RVT U148 ( .A1(N34), .A2(N329), .Y(n152) );
  NAND2X0_RVT U149 ( .A1(N40), .A2(N370), .Y(n151) );
  NAND3X0_RVT U150 ( .A1(n154), .A2(n155), .A3(n156), .Y(n133) );
  NAND2X0_RVT U151 ( .A1(N27), .A2(N370), .Y(n156) );
  NAND2X0_RVT U152 ( .A1(n157), .A2(n158), .Y(n155) );
  NAND2X0_RVT U153 ( .A1(N17), .A2(n159), .Y(n157) );
  NAND2X0_RVT U154 ( .A1(N21), .A2(N329), .Y(n60006) );
  NAND3X0_RVT U155 ( .A1(n160), .A2(n161), .A3(n162), .Y(n141) );
  NAND2X0_RVT U156 ( .A1(N60), .A2(N329), .Y(n161) );
  NAND2X0_RVT U157 ( .A1(N66), .A2(N370), .Y(n160) );
  NAND3X0_RVT U158 ( .A1(n163), .A2(n164), .A3(n165), .Y(n138) );
  NAND2X0_RVT U159 ( .A1(N53), .A2(N370), .Y(n165) );
  NAND2X0_RVT U160 ( .A1(n166), .A2(n167), .Y(n164) );
  NAND2X0_RVT U161 ( .A1(N43), .A2(n159), .Y(n166) );
  NAND2X0_RVT U162 ( .A1(N47), .A2(N329), .Y(n163) );
  NAND2X0_RVT U163 ( .A1(n142), .A2(n146), .Y(n148) );
  NAND3X0_RVT U164 ( .A1(n168), .A2(n169), .A3(n170), .Y(n146) );
  NAND2X0_RVT U165 ( .A1(N92), .A2(N370), .Y(n170) );
  NAND2X0_RVT U166 ( .A1(n171), .A2(n172), .Y(n169) );
  NAND2X0_RVT U167 ( .A1(N82), .A2(n159), .Y(n171) );
  NAND2X0_RVT U168 ( .A1(N86), .A2(N329), .Y(n168) );
  NAND3X0_RVT U169 ( .A1(n173), .A2(n174), .A3(n175), .Y(n142) );
  NAND2X0_RVT U170 ( .A1(N73), .A2(N329), .Y(n174) );
  NAND2X0_RVT U171 ( .A1(N79), .A2(N370), .Y(n173) );
  NAND2X0_RVT U172 ( .A1(n176), .A2(n177), .Y(n145) );
  NAND2X0_RVT U173 ( .A1(N95), .A2(n159), .Y(n177) );
  INVX0_RVT U174 ( .A(N223), .Y(n159) );
  NAND3X0_RVT U175 ( .A1(n178), .A2(n179), .A3(n180), .Y(n149) );
  NAND2X0_RVT U176 ( .A1(N8), .A2(N329), .Y(n179) );
  NAND2X0_RVT U177 ( .A1(N14), .A2(N370), .Y(n178) );
  NAND4X0_RVT U178 ( .A1(n181), .A2(n182), .A3(n183), .A4(n184), .Y(N370) );
  AND4X1_RVT U179 ( .A1(n185), .A2(n186), .A3(n187), .A4(n188), .Y(n184) );
  OR3X1_RVT U180 ( .A1(N115), .A2(n189), .A3(n190), .Y(n188) );
  AND2X1_RVT U181 ( .A1(N329), .A2(n191), .Y(n189) );
  NAND3X0_RVT U182 ( .A1(n192), .A2(n193), .A3(n194), .Y(n187) );
  INVX0_RVT U183 ( .A(N105), .Y(n193) );
  NAND2X0_RVT U184 ( .A1(N329), .A2(n195), .Y(n192) );
  NAND3X0_RVT U185 ( .A1(n196), .A2(n197), .A3(n198), .Y(n186) );
  INVX0_RVT U186 ( .A(N92), .Y(n197) );
  NAND2X0_RVT U187 ( .A1(N329), .A2(n199), .Y(n196) );
  NAND3X0_RVT U188 ( .A1(n200), .A2(n201), .A3(n153), .Y(n185) );
  INVX0_RVT U189 ( .A(N40), .Y(n201) );
  NAND2X0_RVT U190 ( .A1(N329), .A2(n202), .Y(n200) );
  AND3X1_RVT U191 ( .A1(n203), .A2(n204), .A3(n205), .Y(n183) );
  NAND3X0_RVT U192 ( .A1(n206), .A2(n207), .A3(n208), .Y(n205) );
  INVX0_RVT U193 ( .A(N27), .Y(n207) );
  NAND2X0_RVT U194 ( .A1(N329), .A2(n209), .Y(n206) );
  NAND3X0_RVT U195 ( .A1(n210), .A2(n211), .A3(n175), .Y(n204) );
  INVX0_RVT U196 ( .A(N79), .Y(n211) );
  NAND2X0_RVT U197 ( .A1(N329), .A2(n212), .Y(n210) );
  NAND3X0_RVT U198 ( .A1(n213), .A2(n214), .A3(n162), .Y(n203) );
  INVX0_RVT U199 ( .A(N66), .Y(n214) );
  NAND2X0_RVT U200 ( .A1(N329), .A2(n215), .Y(n213) );
  NAND3X0_RVT U201 ( .A1(n216), .A2(n217), .A3(n218), .Y(n182) );
  INVX0_RVT U202 ( .A(N53), .Y(n217) );
  NAND2X0_RVT U203 ( .A1(N329), .A2(n219), .Y(n216) );
  NAND3X0_RVT U204 ( .A1(n220), .A2(n221), .A3(n180), .Y(n181) );
  INVX0_RVT U205 ( .A(N14), .Y(n221) );
  NAND2X0_RVT U206 ( .A1(N329), .A2(n222), .Y(n220) );
  NAND4X0_RVT U207 ( .A1(n202), .A2(n222), .A3(n223), .A4(n224), .Y(N329) );
  AND4X1_RVT U208 ( .A1(n212), .A2(n199), .A3(n195), .A4(n191), .Y(n224) );
  OR2X1_RVT U209 ( .A1(N112), .A2(n190), .Y(n191) );
  NAND2X0_RVT U210 ( .A1(N108), .A2(n225), .Y(n190) );
  NAND2X0_RVT U211 ( .A1(N102), .A2(N223), .Y(n225) );
  AND2X0_RVT U212 ( .A1(n194), .A2(n226), .Y(n60002) );
  INVX0_RVT U213 ( .A(N99), .Y(n226) );
  AND2X1_RVT U214 ( .A1(N95), .A2(n227), .Y(n194) );
  NAND2X0_RVT U215 ( .A1(N223), .A2(n176), .Y(n227) );
  NAND2X0_RVT U216 ( .A1(n198), .A2(n228), .Y(n199) );
  INVX0_RVT U217 ( .A(N86), .Y(n228) );
  AND2X1_RVT U218 ( .A1(N82), .A2(n229), .Y(n60004) );
  NAND2X0_RVT U219 ( .A1(N223), .A2(n172), .Y(n60005) );
  NAND2X0_RVT U220 ( .A1(n175), .A2(n230), .Y(n212) );
  INVX0_RVT U221 ( .A(N73), .Y(n60008) );
  AND2X1_RVT U222 ( .A1(N69), .A2(n231), .Y(n175) );
  NAND2X0_RVT U223 ( .A1(N63), .A2(N223), .Y(n231) );
  AND3X1_RVT U224 ( .A1(n219), .A2(n215), .A3(n209), .Y(n60010) );
  NAND2X0_RVT U225 ( .A1(n208), .A2(n232), .Y(n209) );
  INVX0_RVT U226 ( .A(N21), .Y(n232) );
  AND2X1_RVT U227 ( .A1(N17), .A2(n233), .Y(n208) );
  NAND2X0_RVT U228 ( .A1(N223), .A2(n158), .Y(n233) );
  NAND2X0_RVT U229 ( .A1(n162), .A2(n234), .Y(n215) );
  INVX0_RVT U230 ( .A(N60), .Y(n234) );
  AND2X1_RVT U231 ( .A1(N56), .A2(n235), .Y(n162) );
  NAND2X0_RVT U232 ( .A1(N50), .A2(N223), .Y(n235) );
  NAND2X0_RVT U233 ( .A1(n218), .A2(n236), .Y(n219) );
  INVX0_RVT U234 ( .A(N47), .Y(n236) );
  AND2X1_RVT U235 ( .A1(N43), .A2(n237), .Y(n218) );
  NAND2X0_RVT U236 ( .A1(N223), .A2(n167), .Y(n237) );
  NAND2X0_RVT U237 ( .A1(n180), .A2(n238), .Y(n222) );
  INVX0_RVT U238 ( .A(N8), .Y(n238) );
  AND2X1_RVT U239 ( .A1(N4), .A2(n239), .Y(n180) );
  NAND2X0_RVT U240 ( .A1(N1), .A2(N223), .Y(n239) );
  NAND2X0_RVT U241 ( .A1(n153), .A2(n240), .Y(n202) );
  INVX0_RVT U242 ( .A(N34), .Y(n240) );
  AND2X1_RVT U243 ( .A1(N30), .A2(n241), .Y(n153) );
  NAND2X0_RVT U244 ( .A1(N24), .A2(N223), .Y(n241) );
  NAND4X0_RVT U245 ( .A1(n242), .A2(n172), .A3(n243), .A4(n244), .Y(N223) );
  AND4X1_RVT U246 ( .A1(n245), .A2(n246), .A3(n247), .A4(n248), .Y(n244) );
  NAND2X0_RVT U247 ( .A1(N108), .A2(n249), .Y(n248) );
  INVX0_RVT U248 ( .A(N102), .Y(n249) );
  NAND2X0_RVT U249 ( .A1(N30), .A2(n250), .Y(n60009) );
  INVX0_RVT U250 ( .A(N24), .Y(n250) );
  NAND2X0_RVT U251 ( .A1(N56), .A2(n251), .Y(n246) );
  INVX0_RVT U252 ( .A(N50), .Y(n251) );
  NAND2X0_RVT U253 ( .A1(N69), .A2(n252), .Y(n245) );
  INVX0_RVT U254 ( .A(N63), .Y(n252) );
  AND3X1_RVT U255 ( .A1(n167), .A2(n158), .A3(n176), .Y(n243) );
  NAND2X0_RVT U256 ( .A1(n253), .A2(N95), .Y(n176) );
  INVX0_RVT U257 ( .A(N89), .Y(n253) );
  NAND2X0_RVT U258 ( .A1(n254), .A2(N17), .Y(n158) );
  INVX0_RVT U259 ( .A(N11), .Y(n60003) );
  NAND2X0_RVT U260 ( .A1(n255), .A2(N43), .Y(n167) );
  INVX0_RVT U261 ( .A(N37), .Y(n255) );
  NAND2X0_RVT U262 ( .A1(n256), .A2(N82), .Y(n172) );
  INVX0_RVT U263 ( .A(N76), .Y(n256) );
  NAND2X0_RVT U264 ( .A1(N4), .A2(n257), .Y(n242) );
  INVX0_RVT U265 ( .A(N1), .Y(n257) );
  XOR2X1_RVT U60001 ( .A1(n60001), .A2(1'b1), .Y(n134) );
  XOR2X1_RVT U60002 ( .A1(n60002), .A2(1'b1), .Y(n195) );
  XOR2X1_RVT U60003 ( .A1(n60003), .A2(1'b0), .Y(n254) );
  XOR2X1_RVT U60004 ( .A1(n60004), .A2(1'b0), .Y(n198) );
  XOR2X1_RVT U60005 ( .A1(n60005), .A2(1'b0), .Y(n229) );
  XOR2X1_RVT U60006 ( .A1(n60006), .A2(1'b0), .Y(n154) );
  XOR2X1_RVT U60007 ( .A1(n60007), .A2(1'b0), .Y(n143) );
  XOR2X1_RVT U60008 ( .A1(n60008), .A2(1'b0), .Y(n230) );
  XOR2X1_RVT U60009 ( .A1(n60009), .A2(1'b0), .Y(n247) );
  XOR2X1_RVT U60010 ( .A1(n60010), .A2(1'b0), .Y(n223) );
//new;
endmodule